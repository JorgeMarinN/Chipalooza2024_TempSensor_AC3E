magic
tech sky130A
timestamp 1641587603
<< error_s >>
rect 1466 2536 1506 2576
rect 1426 2496 1466 2536
<< locali >>
rect 2509 3232 2559 3235
rect 2509 3188 2512 3232
rect 2556 3188 2559 3232
rect 2509 3185 2559 3188
<< viali >>
rect 2512 3188 2556 3232
rect 2323 2582 2367 2626
<< metal1 >>
rect 2506 3232 2562 3238
rect 2506 3188 2512 3232
rect 2556 3188 2562 3232
rect 2506 3182 2562 3188
rect 1988 2833 2256 2892
rect 1988 2830 2072 2833
rect 1988 2752 1991 2830
rect 2069 2752 2072 2830
rect 1988 2749 2072 2752
rect 2337 2830 2655 2833
rect 2337 2752 2574 2830
rect 2652 2752 2655 2830
rect 2337 2749 2655 2752
rect 2317 2629 2372 2632
rect 3431 2629 3484 2632
rect 2317 2626 3431 2629
rect 2317 2582 2323 2626
rect 2367 2582 3431 2626
rect 2317 2579 3431 2582
rect 3481 2579 3484 2629
rect 2317 2576 2372 2579
rect 3431 2576 3484 2579
<< via1 >>
rect 1991 2752 2069 2830
rect 2574 2752 2652 2830
rect 3431 2579 3481 2629
<< metal2 >>
rect 1988 2830 2072 2833
rect 1988 2752 1991 2830
rect 2069 2752 2072 2830
rect 1988 2749 2072 2752
rect 2569 2830 2657 2835
rect 2569 2752 2574 2830
rect 2652 2752 2657 2830
rect 2569 2747 2657 2752
rect 3428 2629 3484 2632
rect 3428 2579 3431 2629
rect 3481 2579 3484 2629
rect 3428 2522 3484 2579
<< via2 >>
rect 2574 2752 2652 2830
<< metal3 >>
rect 2570 2830 2873 2833
rect 2570 2752 2574 2830
rect 2652 2752 2792 2830
rect 2870 2752 2873 2830
rect 2570 2749 2873 2752
<< via3 >>
rect 2792 2752 2870 2830
use CAPOSC  CAPOSC_0
timestamp 1641587603
transform 1 0 -1534 0 1 216
box 1534 -216 5016 2653
use INV  INV_0
timestamp 1641587603
transform 1 0 1409 0 1 2683
box 683 -89 1138 540
<< labels >>
flabel space 557 2688 557 2688 0 FreeSans 800 0 0 0 CON_CV
port 1 nsew
flabel space 2247 2896 2247 2896 0 FreeSans 800 0 0 0 VIN
port 2 nsew
flabel via2 2610 2790 2610 2790 0 FreeSans 800 0 0 0 VOUT
port 3 nsew
flabel viali 2517 3196 2517 3196 0 FreeSans 800 0 0 0 VDD
port 4 nsew
flabel metal1 2492 2602 2492 2602 0 FreeSans 800 0 0 0 VSS
port 5 nsew
<< end >>
