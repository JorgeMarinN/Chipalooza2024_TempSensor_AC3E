magic
tech sky130A
magscale 1 2
timestamp 1713593032
<< error_s >>
rect -6020 19649 -5986 23969
rect 682 19649 716 23969
rect 1934 19603 2022 24015
rect 8682 19649 8716 23969
rect 9934 19603 10022 24015
rect 16682 19649 16716 23969
rect -6020 13877 -5986 18197
rect 682 13877 716 18197
rect 1934 13831 2022 18243
rect 8682 13877 8716 18197
rect 9934 13831 10022 18243
rect 16682 13877 16716 18197
rect -6020 8105 -5986 12425
rect 682 8105 716 12425
rect 1934 8059 2022 12471
rect 8682 8105 8716 12425
rect 9934 8059 10022 12471
rect 16682 8105 16716 12425
rect -6020 2333 -5986 6653
rect 682 2333 716 6653
rect 1934 2287 2022 6699
rect 8682 2333 8716 6653
rect 9934 2287 10022 6699
rect 16682 2333 16716 6653
rect -6020 -3439 -5986 881
rect 682 -3439 716 881
rect 1934 -3485 2022 927
rect 8682 -3439 8716 881
rect 9934 -3485 10022 927
rect 16682 -3439 16716 881
rect -8945 -14603 -8909 -14601
rect -8875 -14603 -8839 -14601
rect -7539 -14603 -7447 -14567
rect -6113 -14603 -6021 -14567
rect -4721 -14603 -4685 -14601
rect -4651 -14603 -4615 -14601
rect -8945 -14637 -7503 -14603
rect -7483 -14637 -6077 -14603
rect -6057 -14637 -4615 -14603
rect -8945 -17261 -8909 -14637
rect -8875 -17261 -8839 -14637
rect -7539 -14673 -7447 -14637
rect -6113 -14673 -6021 -14637
rect -7539 -17261 -7447 -17225
rect -6113 -17261 -6021 -17225
rect -4721 -17261 -4685 -14637
rect -4651 -17261 -4615 -14637
rect -8945 -17295 -7503 -17261
rect -7483 -17295 -6077 -17261
rect -6057 -17295 -4615 -17261
rect -8945 -17297 -8909 -17295
rect -8875 -17297 -8839 -17295
rect -7539 -17331 -7447 -17295
rect -6113 -17331 -6021 -17295
rect -4721 -17297 -4685 -17295
rect -4651 -17297 -4615 -17295
<< pdiff >>
rect -6020 -3439 -5986 23969
rect 682 -3439 716 23969
rect 1980 -3439 2014 23969
rect 8682 -3439 8716 23969
rect 9980 -3439 10014 23969
rect 16682 -3439 16716 23969
rect -8909 -14637 -4651 -14603
rect -8909 -17261 -8875 -14637
rect -4685 -17261 -4651 -14637
rect -8909 -17295 -4651 -17261
<< metal1 >>
rect -10661 -1541 -10649 -1529
rect -9846 -4971 -9834 -4959
rect -10051 -7311 -10029 -7289
<< metal2 >>
rect -12332 8816 -7266 9016
rect -10518 1007 -6012 1407
rect -11451 -2121 -11439 -2109
rect -12532 -17430 -7183 -17230
<< metal3 >>
rect -12532 -16042 -9109 -15742
<< metal4 >>
rect -12611 1952 -6666 2152
rect -12611 -10630 -6666 -10430
rect -6866 -14468 -6666 -10630
use ARRAY_RES_HIGH  ARRAY_RES_HIGH_0
timestamp 1713593032
transform 1 0 -8183 0 -1 -15949
box -952 -1481 3758 1481
use ARRAY_RES_ISO  ARRAY_RES_ISO_0
timestamp 1713593032
transform 0 1 -6082 -1 0 17422
box -7073 -1184 21387 24044
use INTERNAL_SDC  INTERNAL_SDC_0
timestamp 1713593032
transform 1 0 -30500 0 1 -11896
box 765 -6413 20802 21798
use vias_gen$16  vias_gen$16_0
timestamp 1713593032
transform 1 0 -12532 0 1 -17430
box 0 0 200 200
use vias_gen$18  vias_gen$18_0
timestamp 1713593032
transform 1 0 -7183 0 1 -17430
box 0 0 800 200
use vias_gen$19  vias_gen$19_0
timestamp 1713593032
transform 1 0 -7183 0 1 -14668
box 0 0 800 200
use vias_gen$21  vias_gen$21_0
timestamp 1713593032
transform 1 0 -12532 0 1 8816
box 0 0 200 200
use vias_gen$24  vias_gen$24_0
timestamp 1713593032
transform 1 0 -6012 0 1 1007
box 0 0 300 400
use vias_gen$25  vias_gen$25_0
timestamp 1713593032
transform 1 0 -6666 0 1 1807
box 0 0 400 400
use vias_gen$26  vias_gen$26_0
timestamp 1713593032
transform 1 0 -10718 0 1 1007
box 0 0 200 400
<< labels >>
flabel metal1 s -10050 -7310 -10030 -7290 2 FreeSans 44 0 0 0 N2_R
port 3 nsew
flabel metal1 s -10660 -1540 -10650 -1530 2 FreeSans 44 0 0 0 VDD
port 1 nsew
flabel metal1 s -12548 8928 -12548 8928 2 FreeSans 44 0 0 0 N3_S
flabel metal1 s -6591 -17363 -6591 -17363 2 FreeSans 44 0 0 0 N3_R
flabel metal1 s -9845 -4970 -9835 -4960 2 FreeSans 44 0 0 0 VSS
port 2 nsew
flabel metal4 s -12179 2044 -12179 2044 2 FreeSans 96 0 0 0 SENS_IN
flabel metal4 s -12102 -10538 -12102 -10538 2 FreeSans 96 0 0 0 REF_IN
flabel metal2 s -11450 -2120 -11440 -2110 2 FreeSans 44 0 0 0 DOUT
port 4 nsew
<< end >>
