magic
tech sky130A
magscale 1 2
timestamp 1713593032
<< metal3 >>
rect -40 1992 2332 2040
rect -40 1928 2248 1992
rect 2312 1928 2332 1992
rect -40 1912 2332 1928
rect -40 1848 2248 1912
rect 2312 1848 2332 1912
rect -40 1832 2332 1848
rect -40 1768 2248 1832
rect 2312 1768 2332 1832
rect -40 1752 2332 1768
rect -40 1688 2248 1752
rect 2312 1688 2332 1752
rect -40 1672 2332 1688
rect -40 1608 2248 1672
rect 2312 1608 2332 1672
rect -40 1592 2332 1608
rect -40 1528 2248 1592
rect 2312 1528 2332 1592
rect -40 1512 2332 1528
rect -40 1448 2248 1512
rect 2312 1448 2332 1512
rect -40 1432 2332 1448
rect -40 1368 2248 1432
rect 2312 1368 2332 1432
rect -40 1352 2332 1368
rect -40 1288 2248 1352
rect 2312 1288 2332 1352
rect -40 1272 2332 1288
rect -40 1208 2248 1272
rect 2312 1208 2332 1272
rect -40 1192 2332 1208
rect -40 1128 2248 1192
rect 2312 1128 2332 1192
rect -40 1112 2332 1128
rect -40 1048 2248 1112
rect 2312 1048 2332 1112
rect -40 1032 2332 1048
rect -40 968 2248 1032
rect 2312 968 2332 1032
rect -40 952 2332 968
rect -40 888 2248 952
rect 2312 888 2332 952
rect -40 872 2332 888
rect -40 808 2248 872
rect 2312 808 2332 872
rect -40 792 2332 808
rect -40 728 2248 792
rect 2312 728 2332 792
rect -40 712 2332 728
rect -40 648 2248 712
rect 2312 648 2332 712
rect -40 632 2332 648
rect -40 568 2248 632
rect 2312 568 2332 632
rect -40 552 2332 568
rect -40 488 2248 552
rect 2312 488 2332 552
rect -40 472 2332 488
rect -40 408 2248 472
rect 2312 408 2332 472
rect -40 392 2332 408
rect -40 328 2248 392
rect 2312 328 2332 392
rect -40 312 2332 328
rect -40 248 2248 312
rect 2312 248 2332 312
rect -40 232 2332 248
rect -40 168 2248 232
rect 2312 168 2332 232
rect -40 152 2332 168
rect -40 88 2248 152
rect 2312 88 2332 152
rect -40 72 2332 88
rect -40 8 2248 72
rect 2312 8 2332 72
rect -40 -40 2332 8
<< via3 >>
rect 2248 1928 2312 1992
rect 2248 1848 2312 1912
rect 2248 1768 2312 1832
rect 2248 1688 2312 1752
rect 2248 1608 2312 1672
rect 2248 1528 2312 1592
rect 2248 1448 2312 1512
rect 2248 1368 2312 1432
rect 2248 1288 2312 1352
rect 2248 1208 2312 1272
rect 2248 1128 2312 1192
rect 2248 1048 2312 1112
rect 2248 968 2312 1032
rect 2248 888 2312 952
rect 2248 808 2312 872
rect 2248 728 2312 792
rect 2248 648 2312 712
rect 2248 568 2312 632
rect 2248 488 2312 552
rect 2248 408 2312 472
rect 2248 328 2312 392
rect 2248 248 2312 312
rect 2248 168 2312 232
rect 2248 88 2312 152
rect 2248 8 2312 72
<< mimcap >>
rect 0 1952 2000 2000
rect 0 48 48 1952
rect 1952 48 2000 1952
rect 0 0 2000 48
<< mimcapcontact >>
rect 48 48 1952 1952
<< metal4 >>
rect 2232 1992 2328 2028
rect 39 1952 1961 1961
rect 39 48 48 1952
rect 1952 48 1961 1952
rect 39 39 1961 48
rect 2232 1928 2248 1992
rect 2312 1928 2328 1992
rect 2232 1912 2328 1928
rect 2232 1848 2248 1912
rect 2312 1848 2328 1912
rect 2232 1832 2328 1848
rect 2232 1768 2248 1832
rect 2312 1768 2328 1832
rect 2232 1752 2328 1768
rect 2232 1688 2248 1752
rect 2312 1688 2328 1752
rect 2232 1672 2328 1688
rect 2232 1608 2248 1672
rect 2312 1608 2328 1672
rect 2232 1592 2328 1608
rect 2232 1528 2248 1592
rect 2312 1528 2328 1592
rect 2232 1512 2328 1528
rect 2232 1448 2248 1512
rect 2312 1448 2328 1512
rect 2232 1432 2328 1448
rect 2232 1368 2248 1432
rect 2312 1368 2328 1432
rect 2232 1352 2328 1368
rect 2232 1288 2248 1352
rect 2312 1288 2328 1352
rect 2232 1272 2328 1288
rect 2232 1208 2248 1272
rect 2312 1208 2328 1272
rect 2232 1192 2328 1208
rect 2232 1128 2248 1192
rect 2312 1128 2328 1192
rect 2232 1112 2328 1128
rect 2232 1048 2248 1112
rect 2312 1048 2328 1112
rect 2232 1032 2328 1048
rect 2232 968 2248 1032
rect 2312 968 2328 1032
rect 2232 952 2328 968
rect 2232 888 2248 952
rect 2312 888 2328 952
rect 2232 872 2328 888
rect 2232 808 2248 872
rect 2312 808 2328 872
rect 2232 792 2328 808
rect 2232 728 2248 792
rect 2312 728 2328 792
rect 2232 712 2328 728
rect 2232 648 2248 712
rect 2312 648 2328 712
rect 2232 632 2328 648
rect 2232 568 2248 632
rect 2312 568 2328 632
rect 2232 552 2328 568
rect 2232 488 2248 552
rect 2312 488 2328 552
rect 2232 472 2328 488
rect 2232 408 2248 472
rect 2312 408 2328 472
rect 2232 392 2328 408
rect 2232 328 2248 392
rect 2312 328 2328 392
rect 2232 312 2328 328
rect 2232 248 2248 312
rect 2312 248 2328 312
rect 2232 232 2328 248
rect 2232 168 2248 232
rect 2312 168 2328 232
rect 2232 152 2328 168
rect 2232 88 2248 152
rect 2312 88 2328 152
rect 2232 72 2328 88
rect 2232 8 2248 72
rect 2312 8 2328 72
rect 2232 -28 2328 8
<< end >>
