magic
tech sky130A
timestamp 1713591521
<< metal1 >>
rect 0 193 150 200
rect 0 7 14 193
rect 136 7 150 193
rect 0 0 150 7
<< via1 >>
rect 14 7 136 193
<< metal2 >>
rect 0 193 150 200
rect 0 7 14 193
rect 136 7 150 193
rect 0 0 150 7
<< end >>
