magic
tech sky130A
magscale 1 2
timestamp 1713591521
<< poly >>
rect 0 151 66 200
rect 0 117 16 151
rect 50 117 66 151
rect 0 83 66 117
rect 0 49 16 83
rect 50 49 66 83
rect 0 0 66 49
<< polycont >>
rect 16 117 50 151
rect 16 49 50 83
<< locali >>
rect 0 153 66 200
rect 0 117 16 153
rect 50 117 66 153
rect 0 83 66 117
rect 0 47 16 83
rect 50 47 66 83
rect 0 0 66 47
<< viali >>
rect 16 151 50 153
rect 16 119 50 151
rect 16 49 50 81
rect 16 47 50 49
<< metal1 >>
rect 0 153 66 200
rect 0 119 16 153
rect 50 119 66 153
rect 0 81 66 119
rect 0 47 16 81
rect 50 47 66 81
rect 0 0 66 47
<< end >>
