magic
tech sky130A
magscale 1 2
timestamp 1713591521
<< error_s >>
rect -6001 19628 -5967 23948
rect 701 19628 735 23948
rect 1999 19628 2033 23948
rect 8701 19628 8735 23948
rect 9999 19628 10033 23948
rect 16701 19628 16735 23948
rect -6001 13856 -5967 18176
rect 701 13856 735 18176
rect 1999 13856 2033 18176
rect 8701 13856 8735 18176
rect 9999 13856 10033 18176
rect 16701 13856 16735 18176
rect -14853 9861 -14797 9881
rect -14773 9861 -14717 9881
rect -14885 9805 -14853 9861
rect -14797 9805 -14773 9861
rect -14717 9805 -14685 9861
rect -14853 9621 -14797 9805
rect -14773 9621 -14717 9805
rect -6001 8084 -5967 12404
rect 701 8084 735 12404
rect 1999 8084 2033 12404
rect 8701 8084 8735 12404
rect 9999 8084 10033 12404
rect 16701 8084 16735 12404
rect -6001 2312 -5967 6632
rect 701 2312 735 6632
rect 1999 2312 2033 6632
rect 8701 2312 8735 6632
rect 9999 2312 10033 6632
rect 16701 2312 16735 6632
rect -6001 -3460 -5967 860
rect 701 -3460 735 860
rect 1999 -3460 2033 860
rect 8701 -3460 8735 860
rect 9999 -3460 10033 860
rect 16701 -3460 16735 860
rect -8926 -14624 -8890 -14622
rect -8856 -14624 -8820 -14622
rect -7520 -14624 -7428 -14588
rect -6094 -14624 -6002 -14588
rect -4702 -14624 -4666 -14622
rect -4632 -14624 -4596 -14622
rect -8926 -14658 -7484 -14624
rect -7464 -14658 -6058 -14624
rect -6038 -14658 -4596 -14624
rect -8926 -17282 -8890 -14658
rect -8856 -17282 -8820 -14658
rect -7520 -14694 -7428 -14658
rect -6094 -14694 -6002 -14658
rect -7520 -17282 -7428 -17246
rect -6094 -17282 -6002 -17246
rect -4702 -17282 -4666 -14658
rect -4632 -17282 -4596 -14658
rect -8926 -17316 -7484 -17282
rect -7464 -17316 -6058 -17282
rect -6038 -17316 -4596 -17282
rect -8926 -17318 -8890 -17316
rect -8856 -17318 -8820 -17316
rect -7520 -17352 -7428 -17316
rect -6094 -17352 -6002 -17316
rect -4702 -17318 -4666 -17316
rect -4632 -17318 -4596 -17316
rect -14853 -18254 -14797 -18070
rect -14773 -18254 -14717 -18070
rect -14885 -18310 -14853 -18254
rect -14797 -18310 -14773 -18254
rect -14717 -18310 -14685 -18254
rect -14853 -18330 -14797 -18310
rect -14773 -18330 -14717 -18310
<< dnwell >>
rect -30116 -18730 18381 24874
<< nwell >>
rect -30196 24668 18461 24954
rect -30196 -18524 -29910 24668
rect 18175 -18524 18461 24668
rect -30196 -18810 18461 -18524
<< nsubdiff >>
rect -29910 24848 -29750 24874
rect -29910 24808 -29880 24848
rect -29840 24808 -29806 24848
rect -29766 24808 -29750 24848
rect -29910 24774 -29750 24808
rect -29910 24734 -29880 24774
rect -29840 24734 -29806 24774
rect -29766 24734 -29750 24774
rect -29910 24704 -29750 24734
rect -27910 24848 -27750 24874
rect -27910 24808 -27880 24848
rect -27840 24808 -27806 24848
rect -27766 24808 -27750 24848
rect -27910 24774 -27750 24808
rect -27910 24734 -27880 24774
rect -27840 24734 -27806 24774
rect -27766 24734 -27750 24774
rect -27910 24704 -27750 24734
rect -25910 24848 -25750 24874
rect -25910 24808 -25880 24848
rect -25840 24808 -25806 24848
rect -25766 24808 -25750 24848
rect -25910 24774 -25750 24808
rect -25910 24734 -25880 24774
rect -25840 24734 -25806 24774
rect -25766 24734 -25750 24774
rect -25910 24704 -25750 24734
rect -23910 24848 -23750 24874
rect -23910 24808 -23880 24848
rect -23840 24808 -23806 24848
rect -23766 24808 -23750 24848
rect -23910 24774 -23750 24808
rect -23910 24734 -23880 24774
rect -23840 24734 -23806 24774
rect -23766 24734 -23750 24774
rect -23910 24704 -23750 24734
rect -21910 24848 -21750 24874
rect -21910 24808 -21880 24848
rect -21840 24808 -21806 24848
rect -21766 24808 -21750 24848
rect -21910 24774 -21750 24808
rect -21910 24734 -21880 24774
rect -21840 24734 -21806 24774
rect -21766 24734 -21750 24774
rect -21910 24704 -21750 24734
rect -19910 24848 -19750 24874
rect -19910 24808 -19880 24848
rect -19840 24808 -19806 24848
rect -19766 24808 -19750 24848
rect -19910 24774 -19750 24808
rect -19910 24734 -19880 24774
rect -19840 24734 -19806 24774
rect -19766 24734 -19750 24774
rect -19910 24704 -19750 24734
rect -17910 24848 -17750 24874
rect -17910 24808 -17880 24848
rect -17840 24808 -17806 24848
rect -17766 24808 -17750 24848
rect -17910 24774 -17750 24808
rect -17910 24734 -17880 24774
rect -17840 24734 -17806 24774
rect -17766 24734 -17750 24774
rect -17910 24704 -17750 24734
rect -15910 24848 -15750 24874
rect -15910 24808 -15880 24848
rect -15840 24808 -15806 24848
rect -15766 24808 -15750 24848
rect -15910 24774 -15750 24808
rect -15910 24734 -15880 24774
rect -15840 24734 -15806 24774
rect -15766 24734 -15750 24774
rect -15910 24704 -15750 24734
rect -13910 24848 -13750 24874
rect -13910 24808 -13880 24848
rect -13840 24808 -13806 24848
rect -13766 24808 -13750 24848
rect -13910 24774 -13750 24808
rect -13910 24734 -13880 24774
rect -13840 24734 -13806 24774
rect -13766 24734 -13750 24774
rect -13910 24704 -13750 24734
rect -11910 24848 -11750 24874
rect -11910 24808 -11880 24848
rect -11840 24808 -11806 24848
rect -11766 24808 -11750 24848
rect -11910 24774 -11750 24808
rect -11910 24734 -11880 24774
rect -11840 24734 -11806 24774
rect -11766 24734 -11750 24774
rect -11910 24704 -11750 24734
rect -9910 24848 -9750 24874
rect -9910 24808 -9880 24848
rect -9840 24808 -9806 24848
rect -9766 24808 -9750 24848
rect -9910 24774 -9750 24808
rect -9910 24734 -9880 24774
rect -9840 24734 -9806 24774
rect -9766 24734 -9750 24774
rect -9910 24704 -9750 24734
rect -7910 24848 -7750 24874
rect -7910 24808 -7880 24848
rect -7840 24808 -7806 24848
rect -7766 24808 -7750 24848
rect -7910 24774 -7750 24808
rect -7910 24734 -7880 24774
rect -7840 24734 -7806 24774
rect -7766 24734 -7750 24774
rect -7910 24704 -7750 24734
rect -5910 24848 -5750 24874
rect -5910 24808 -5880 24848
rect -5840 24808 -5806 24848
rect -5766 24808 -5750 24848
rect -5910 24774 -5750 24808
rect -5910 24734 -5880 24774
rect -5840 24734 -5806 24774
rect -5766 24734 -5750 24774
rect -5910 24704 -5750 24734
rect -3910 24848 -3750 24874
rect -3910 24808 -3880 24848
rect -3840 24808 -3806 24848
rect -3766 24808 -3750 24848
rect -3910 24774 -3750 24808
rect -3910 24734 -3880 24774
rect -3840 24734 -3806 24774
rect -3766 24734 -3750 24774
rect -3910 24704 -3750 24734
rect -1910 24848 -1750 24874
rect -1910 24808 -1880 24848
rect -1840 24808 -1806 24848
rect -1766 24808 -1750 24848
rect -1910 24774 -1750 24808
rect -1910 24734 -1880 24774
rect -1840 24734 -1806 24774
rect -1766 24734 -1750 24774
rect -1910 24704 -1750 24734
rect 90 24848 250 24874
rect 90 24808 120 24848
rect 160 24808 194 24848
rect 234 24808 250 24848
rect 90 24774 250 24808
rect 90 24734 120 24774
rect 160 24734 194 24774
rect 234 24734 250 24774
rect 90 24704 250 24734
rect 2090 24848 2250 24874
rect 2090 24808 2120 24848
rect 2160 24808 2194 24848
rect 2234 24808 2250 24848
rect 2090 24774 2250 24808
rect 2090 24734 2120 24774
rect 2160 24734 2194 24774
rect 2234 24734 2250 24774
rect 2090 24704 2250 24734
rect 4090 24848 4250 24874
rect 4090 24808 4120 24848
rect 4160 24808 4194 24848
rect 4234 24808 4250 24848
rect 4090 24774 4250 24808
rect 4090 24734 4120 24774
rect 4160 24734 4194 24774
rect 4234 24734 4250 24774
rect 4090 24704 4250 24734
rect 6090 24848 6250 24874
rect 6090 24808 6120 24848
rect 6160 24808 6194 24848
rect 6234 24808 6250 24848
rect 6090 24774 6250 24808
rect 6090 24734 6120 24774
rect 6160 24734 6194 24774
rect 6234 24734 6250 24774
rect 6090 24704 6250 24734
rect 8090 24848 8250 24874
rect 8090 24808 8120 24848
rect 8160 24808 8194 24848
rect 8234 24808 8250 24848
rect 8090 24774 8250 24808
rect 8090 24734 8120 24774
rect 8160 24734 8194 24774
rect 8234 24734 8250 24774
rect 8090 24704 8250 24734
rect 10090 24848 10250 24874
rect 10090 24808 10120 24848
rect 10160 24808 10194 24848
rect 10234 24808 10250 24848
rect 10090 24774 10250 24808
rect 10090 24734 10120 24774
rect 10160 24734 10194 24774
rect 10234 24734 10250 24774
rect 10090 24704 10250 24734
rect 12090 24848 12250 24874
rect 12090 24808 12120 24848
rect 12160 24808 12194 24848
rect 12234 24808 12250 24848
rect 12090 24774 12250 24808
rect 12090 24734 12120 24774
rect 12160 24734 12194 24774
rect 12234 24734 12250 24774
rect 12090 24704 12250 24734
rect 14090 24848 14250 24874
rect 14090 24808 14120 24848
rect 14160 24808 14194 24848
rect 14234 24808 14250 24848
rect 14090 24774 14250 24808
rect 14090 24734 14120 24774
rect 14160 24734 14194 24774
rect 14234 24734 14250 24774
rect 14090 24704 14250 24734
rect 16090 24848 16250 24874
rect 16090 24808 16120 24848
rect 16160 24808 16194 24848
rect 16234 24808 16250 24848
rect 16090 24774 16250 24808
rect 16090 24734 16120 24774
rect 16160 24734 16194 24774
rect 16234 24734 16250 24774
rect 16090 24704 16250 24734
rect 18090 24848 18250 24874
rect 18090 24808 18120 24848
rect 18160 24808 18194 24848
rect 18234 24808 18250 24848
rect 18090 24774 18250 24808
rect 18090 24734 18120 24774
rect 18160 24734 18194 24774
rect 18234 24734 18250 24774
rect 18090 24704 18250 24734
rect 18220 24120 18380 24146
rect 18220 24080 18250 24120
rect 18290 24080 18324 24120
rect 18364 24080 18380 24120
rect 18220 24046 18380 24080
rect 18220 24006 18250 24046
rect 18290 24006 18324 24046
rect 18364 24006 18380 24046
rect 18220 23976 18380 24006
rect -30116 23630 -29956 23656
rect -30116 23590 -30086 23630
rect -30046 23590 -30012 23630
rect -29972 23590 -29956 23630
rect -30116 23556 -29956 23590
rect -30116 23516 -30086 23556
rect -30046 23516 -30012 23556
rect -29972 23516 -29956 23556
rect -30116 23486 -29956 23516
rect 18220 22120 18380 22146
rect 18220 22080 18250 22120
rect 18290 22080 18324 22120
rect 18364 22080 18380 22120
rect 18220 22046 18380 22080
rect 18220 22006 18250 22046
rect 18290 22006 18324 22046
rect 18364 22006 18380 22046
rect 18220 21976 18380 22006
rect -30116 21630 -29956 21656
rect -30116 21590 -30086 21630
rect -30046 21590 -30012 21630
rect -29972 21590 -29956 21630
rect -30116 21556 -29956 21590
rect -30116 21516 -30086 21556
rect -30046 21516 -30012 21556
rect -29972 21516 -29956 21556
rect -30116 21486 -29956 21516
rect 18220 20120 18380 20146
rect 18220 20080 18250 20120
rect 18290 20080 18324 20120
rect 18364 20080 18380 20120
rect 18220 20046 18380 20080
rect 18220 20006 18250 20046
rect 18290 20006 18324 20046
rect 18364 20006 18380 20046
rect 18220 19976 18380 20006
rect -30116 19630 -29956 19656
rect -30116 19590 -30086 19630
rect -30046 19590 -30012 19630
rect -29972 19590 -29956 19630
rect -30116 19556 -29956 19590
rect -30116 19516 -30086 19556
rect -30046 19516 -30012 19556
rect -29972 19516 -29956 19556
rect -30116 19486 -29956 19516
rect 18220 18120 18380 18146
rect 18220 18080 18250 18120
rect 18290 18080 18324 18120
rect 18364 18080 18380 18120
rect 18220 18046 18380 18080
rect 18220 18006 18250 18046
rect 18290 18006 18324 18046
rect 18364 18006 18380 18046
rect 18220 17976 18380 18006
rect -30116 17630 -29956 17656
rect -30116 17590 -30086 17630
rect -30046 17590 -30012 17630
rect -29972 17590 -29956 17630
rect -30116 17556 -29956 17590
rect -30116 17516 -30086 17556
rect -30046 17516 -30012 17556
rect -29972 17516 -29956 17556
rect -30116 17486 -29956 17516
rect 18220 16120 18380 16146
rect 18220 16080 18250 16120
rect 18290 16080 18324 16120
rect 18364 16080 18380 16120
rect 18220 16046 18380 16080
rect 18220 16006 18250 16046
rect 18290 16006 18324 16046
rect 18364 16006 18380 16046
rect 18220 15976 18380 16006
rect -30116 15630 -29956 15656
rect -30116 15590 -30086 15630
rect -30046 15590 -30012 15630
rect -29972 15590 -29956 15630
rect -30116 15556 -29956 15590
rect -30116 15516 -30086 15556
rect -30046 15516 -30012 15556
rect -29972 15516 -29956 15556
rect -30116 15486 -29956 15516
rect 18220 14120 18380 14146
rect 18220 14080 18250 14120
rect 18290 14080 18324 14120
rect 18364 14080 18380 14120
rect 18220 14046 18380 14080
rect 18220 14006 18250 14046
rect 18290 14006 18324 14046
rect 18364 14006 18380 14046
rect 18220 13976 18380 14006
rect -30116 13630 -29956 13656
rect -30116 13590 -30086 13630
rect -30046 13590 -30012 13630
rect -29972 13590 -29956 13630
rect -30116 13556 -29956 13590
rect -30116 13516 -30086 13556
rect -30046 13516 -30012 13556
rect -29972 13516 -29956 13556
rect -30116 13486 -29956 13516
rect 18220 12120 18380 12146
rect 18220 12080 18250 12120
rect 18290 12080 18324 12120
rect 18364 12080 18380 12120
rect 18220 12046 18380 12080
rect 18220 12006 18250 12046
rect 18290 12006 18324 12046
rect 18364 12006 18380 12046
rect 18220 11976 18380 12006
rect -30116 11630 -29956 11656
rect -30116 11590 -30086 11630
rect -30046 11590 -30012 11630
rect -29972 11590 -29956 11630
rect -30116 11556 -29956 11590
rect -30116 11516 -30086 11556
rect -30046 11516 -30012 11556
rect -29972 11516 -29956 11556
rect -30116 11486 -29956 11516
rect 18220 10120 18380 10146
rect 18220 10080 18250 10120
rect 18290 10080 18324 10120
rect 18364 10080 18380 10120
rect 18220 10046 18380 10080
rect 18220 10006 18250 10046
rect 18290 10006 18324 10046
rect 18364 10006 18380 10046
rect 18220 9976 18380 10006
rect -30116 9630 -29956 9656
rect -30116 9590 -30086 9630
rect -30046 9590 -30012 9630
rect -29972 9590 -29956 9630
rect -30116 9556 -29956 9590
rect -30116 9516 -30086 9556
rect -30046 9516 -30012 9556
rect -29972 9516 -29956 9556
rect -30116 9486 -29956 9516
rect 18220 8120 18380 8146
rect 18220 8080 18250 8120
rect 18290 8080 18324 8120
rect 18364 8080 18380 8120
rect 18220 8046 18380 8080
rect 18220 8006 18250 8046
rect 18290 8006 18324 8046
rect 18364 8006 18380 8046
rect 18220 7976 18380 8006
rect -30116 7630 -29956 7656
rect -30116 7590 -30086 7630
rect -30046 7590 -30012 7630
rect -29972 7590 -29956 7630
rect -30116 7556 -29956 7590
rect -30116 7516 -30086 7556
rect -30046 7516 -30012 7556
rect -29972 7516 -29956 7556
rect -30116 7486 -29956 7516
rect 18220 6120 18380 6146
rect 18220 6080 18250 6120
rect 18290 6080 18324 6120
rect 18364 6080 18380 6120
rect 18220 6046 18380 6080
rect 18220 6006 18250 6046
rect 18290 6006 18324 6046
rect 18364 6006 18380 6046
rect 18220 5976 18380 6006
rect -30116 5630 -29956 5656
rect -30116 5590 -30086 5630
rect -30046 5590 -30012 5630
rect -29972 5590 -29956 5630
rect -30116 5556 -29956 5590
rect -30116 5516 -30086 5556
rect -30046 5516 -30012 5556
rect -29972 5516 -29956 5556
rect -30116 5486 -29956 5516
rect 18220 4120 18380 4146
rect 18220 4080 18250 4120
rect 18290 4080 18324 4120
rect 18364 4080 18380 4120
rect 18220 4046 18380 4080
rect 18220 4006 18250 4046
rect 18290 4006 18324 4046
rect 18364 4006 18380 4046
rect 18220 3976 18380 4006
rect -30116 3630 -29956 3656
rect -30116 3590 -30086 3630
rect -30046 3590 -30012 3630
rect -29972 3590 -29956 3630
rect -30116 3556 -29956 3590
rect -30116 3516 -30086 3556
rect -30046 3516 -30012 3556
rect -29972 3516 -29956 3556
rect -30116 3486 -29956 3516
rect 18220 2120 18380 2146
rect 18220 2080 18250 2120
rect 18290 2080 18324 2120
rect 18364 2080 18380 2120
rect 18220 2046 18380 2080
rect 18220 2006 18250 2046
rect 18290 2006 18324 2046
rect 18364 2006 18380 2046
rect 18220 1976 18380 2006
rect -30116 1630 -29956 1656
rect -30116 1590 -30086 1630
rect -30046 1590 -30012 1630
rect -29972 1590 -29956 1630
rect -30116 1556 -29956 1590
rect -30116 1516 -30086 1556
rect -30046 1516 -30012 1556
rect -29972 1516 -29956 1556
rect -30116 1486 -29956 1516
rect 18220 120 18380 146
rect 18220 80 18250 120
rect 18290 80 18324 120
rect 18364 80 18380 120
rect 18220 46 18380 80
rect 18220 6 18250 46
rect 18290 6 18324 46
rect 18364 6 18380 46
rect 18220 -24 18380 6
rect -30116 -370 -29956 -344
rect -30116 -410 -30086 -370
rect -30046 -410 -30012 -370
rect -29972 -410 -29956 -370
rect -30116 -444 -29956 -410
rect -30116 -484 -30086 -444
rect -30046 -484 -30012 -444
rect -29972 -484 -29956 -444
rect -30116 -514 -29956 -484
rect 18220 -1880 18380 -1854
rect 18220 -1920 18250 -1880
rect 18290 -1920 18324 -1880
rect 18364 -1920 18380 -1880
rect 18220 -1954 18380 -1920
rect 18220 -1994 18250 -1954
rect 18290 -1994 18324 -1954
rect 18364 -1994 18380 -1954
rect 18220 -2024 18380 -1994
rect -30116 -2370 -29956 -2344
rect -30116 -2410 -30086 -2370
rect -30046 -2410 -30012 -2370
rect -29972 -2410 -29956 -2370
rect -30116 -2444 -29956 -2410
rect -30116 -2484 -30086 -2444
rect -30046 -2484 -30012 -2444
rect -29972 -2484 -29956 -2444
rect -30116 -2514 -29956 -2484
rect 18220 -3880 18380 -3854
rect 18220 -3920 18250 -3880
rect 18290 -3920 18324 -3880
rect 18364 -3920 18380 -3880
rect 18220 -3954 18380 -3920
rect 18220 -3994 18250 -3954
rect 18290 -3994 18324 -3954
rect 18364 -3994 18380 -3954
rect 18220 -4024 18380 -3994
rect -30116 -4370 -29956 -4344
rect -30116 -4410 -30086 -4370
rect -30046 -4410 -30012 -4370
rect -29972 -4410 -29956 -4370
rect -30116 -4444 -29956 -4410
rect -30116 -4484 -30086 -4444
rect -30046 -4484 -30012 -4444
rect -29972 -4484 -29956 -4444
rect -30116 -4514 -29956 -4484
rect 18220 -5880 18380 -5854
rect 18220 -5920 18250 -5880
rect 18290 -5920 18324 -5880
rect 18364 -5920 18380 -5880
rect 18220 -5954 18380 -5920
rect 18220 -5994 18250 -5954
rect 18290 -5994 18324 -5954
rect 18364 -5994 18380 -5954
rect 18220 -6024 18380 -5994
rect -30116 -6370 -29956 -6344
rect -30116 -6410 -30086 -6370
rect -30046 -6410 -30012 -6370
rect -29972 -6410 -29956 -6370
rect -30116 -6444 -29956 -6410
rect -30116 -6484 -30086 -6444
rect -30046 -6484 -30012 -6444
rect -29972 -6484 -29956 -6444
rect -30116 -6514 -29956 -6484
rect 18220 -7880 18380 -7854
rect 18220 -7920 18250 -7880
rect 18290 -7920 18324 -7880
rect 18364 -7920 18380 -7880
rect 18220 -7954 18380 -7920
rect 18220 -7994 18250 -7954
rect 18290 -7994 18324 -7954
rect 18364 -7994 18380 -7954
rect 18220 -8024 18380 -7994
rect -30116 -8370 -29956 -8344
rect -30116 -8410 -30086 -8370
rect -30046 -8410 -30012 -8370
rect -29972 -8410 -29956 -8370
rect -30116 -8444 -29956 -8410
rect -30116 -8484 -30086 -8444
rect -30046 -8484 -30012 -8444
rect -29972 -8484 -29956 -8444
rect -30116 -8514 -29956 -8484
rect 18220 -9880 18380 -9854
rect 18220 -9920 18250 -9880
rect 18290 -9920 18324 -9880
rect 18364 -9920 18380 -9880
rect 18220 -9954 18380 -9920
rect 18220 -9994 18250 -9954
rect 18290 -9994 18324 -9954
rect 18364 -9994 18380 -9954
rect 18220 -10024 18380 -9994
rect -30116 -10370 -29956 -10344
rect -30116 -10410 -30086 -10370
rect -30046 -10410 -30012 -10370
rect -29972 -10410 -29956 -10370
rect -30116 -10444 -29956 -10410
rect -30116 -10484 -30086 -10444
rect -30046 -10484 -30012 -10444
rect -29972 -10484 -29956 -10444
rect -30116 -10514 -29956 -10484
rect 18220 -11880 18380 -11854
rect 18220 -11920 18250 -11880
rect 18290 -11920 18324 -11880
rect 18364 -11920 18380 -11880
rect 18220 -11954 18380 -11920
rect 18220 -11994 18250 -11954
rect 18290 -11994 18324 -11954
rect 18364 -11994 18380 -11954
rect 18220 -12024 18380 -11994
rect -30116 -12370 -29956 -12344
rect -30116 -12410 -30086 -12370
rect -30046 -12410 -30012 -12370
rect -29972 -12410 -29956 -12370
rect -30116 -12444 -29956 -12410
rect -30116 -12484 -30086 -12444
rect -30046 -12484 -30012 -12444
rect -29972 -12484 -29956 -12444
rect -30116 -12514 -29956 -12484
rect 18220 -13880 18380 -13854
rect 18220 -13920 18250 -13880
rect 18290 -13920 18324 -13880
rect 18364 -13920 18380 -13880
rect 18220 -13954 18380 -13920
rect 18220 -13994 18250 -13954
rect 18290 -13994 18324 -13954
rect 18364 -13994 18380 -13954
rect 18220 -14024 18380 -13994
rect -30116 -14370 -29956 -14344
rect -30116 -14410 -30086 -14370
rect -30046 -14410 -30012 -14370
rect -29972 -14410 -29956 -14370
rect -30116 -14444 -29956 -14410
rect -30116 -14484 -30086 -14444
rect -30046 -14484 -30012 -14444
rect -29972 -14484 -29956 -14444
rect -30116 -14514 -29956 -14484
rect 18220 -15880 18380 -15854
rect 18220 -15920 18250 -15880
rect 18290 -15920 18324 -15880
rect 18364 -15920 18380 -15880
rect 18220 -15954 18380 -15920
rect 18220 -15994 18250 -15954
rect 18290 -15994 18324 -15954
rect 18364 -15994 18380 -15954
rect 18220 -16024 18380 -15994
rect -30116 -16370 -29956 -16344
rect -30116 -16410 -30086 -16370
rect -30046 -16410 -30012 -16370
rect -29972 -16410 -29956 -16370
rect -30116 -16444 -29956 -16410
rect -30116 -16484 -30086 -16444
rect -30046 -16484 -30012 -16444
rect -29972 -16484 -29956 -16444
rect -30116 -16514 -29956 -16484
rect 18220 -17880 18380 -17854
rect 18220 -17920 18250 -17880
rect 18290 -17920 18324 -17880
rect 18364 -17920 18380 -17880
rect 18220 -17954 18380 -17920
rect 18220 -17994 18250 -17954
rect 18290 -17994 18324 -17954
rect 18364 -17994 18380 -17954
rect 18220 -18024 18380 -17994
rect -30116 -18370 -29956 -18344
rect -30116 -18410 -30086 -18370
rect -30046 -18410 -30012 -18370
rect -29972 -18410 -29956 -18370
rect -30116 -18444 -29956 -18410
rect -30116 -18484 -30086 -18444
rect -30046 -18484 -30012 -18444
rect -29972 -18484 -29956 -18444
rect -30116 -18514 -29956 -18484
rect -28930 -18586 -28770 -18560
rect -28930 -18626 -28900 -18586
rect -28860 -18626 -28826 -18586
rect -28786 -18626 -28770 -18586
rect -28930 -18660 -28770 -18626
rect -28930 -18700 -28900 -18660
rect -28860 -18700 -28826 -18660
rect -28786 -18700 -28770 -18660
rect -28930 -18730 -28770 -18700
rect -26930 -18586 -26770 -18560
rect -26930 -18626 -26900 -18586
rect -26860 -18626 -26826 -18586
rect -26786 -18626 -26770 -18586
rect -26930 -18660 -26770 -18626
rect -26930 -18700 -26900 -18660
rect -26860 -18700 -26826 -18660
rect -26786 -18700 -26770 -18660
rect -26930 -18730 -26770 -18700
rect -24930 -18586 -24770 -18560
rect -24930 -18626 -24900 -18586
rect -24860 -18626 -24826 -18586
rect -24786 -18626 -24770 -18586
rect -24930 -18660 -24770 -18626
rect -24930 -18700 -24900 -18660
rect -24860 -18700 -24826 -18660
rect -24786 -18700 -24770 -18660
rect -24930 -18730 -24770 -18700
rect -22930 -18586 -22770 -18560
rect -22930 -18626 -22900 -18586
rect -22860 -18626 -22826 -18586
rect -22786 -18626 -22770 -18586
rect -22930 -18660 -22770 -18626
rect -22930 -18700 -22900 -18660
rect -22860 -18700 -22826 -18660
rect -22786 -18700 -22770 -18660
rect -22930 -18730 -22770 -18700
rect -20930 -18586 -20770 -18560
rect -20930 -18626 -20900 -18586
rect -20860 -18626 -20826 -18586
rect -20786 -18626 -20770 -18586
rect -20930 -18660 -20770 -18626
rect -20930 -18700 -20900 -18660
rect -20860 -18700 -20826 -18660
rect -20786 -18700 -20770 -18660
rect -20930 -18730 -20770 -18700
rect -18930 -18586 -18770 -18560
rect -18930 -18626 -18900 -18586
rect -18860 -18626 -18826 -18586
rect -18786 -18626 -18770 -18586
rect -18930 -18660 -18770 -18626
rect -18930 -18700 -18900 -18660
rect -18860 -18700 -18826 -18660
rect -18786 -18700 -18770 -18660
rect -18930 -18730 -18770 -18700
rect -16930 -18586 -16770 -18560
rect -16930 -18626 -16900 -18586
rect -16860 -18626 -16826 -18586
rect -16786 -18626 -16770 -18586
rect -16930 -18660 -16770 -18626
rect -16930 -18700 -16900 -18660
rect -16860 -18700 -16826 -18660
rect -16786 -18700 -16770 -18660
rect -16930 -18730 -16770 -18700
rect -14930 -18586 -14770 -18560
rect -14930 -18626 -14900 -18586
rect -14860 -18626 -14826 -18586
rect -14786 -18626 -14770 -18586
rect -14930 -18660 -14770 -18626
rect -14930 -18700 -14900 -18660
rect -14860 -18700 -14826 -18660
rect -14786 -18700 -14770 -18660
rect -14930 -18730 -14770 -18700
rect -12930 -18586 -12770 -18560
rect -12930 -18626 -12900 -18586
rect -12860 -18626 -12826 -18586
rect -12786 -18626 -12770 -18586
rect -12930 -18660 -12770 -18626
rect -12930 -18700 -12900 -18660
rect -12860 -18700 -12826 -18660
rect -12786 -18700 -12770 -18660
rect -12930 -18730 -12770 -18700
rect -10930 -18586 -10770 -18560
rect -10930 -18626 -10900 -18586
rect -10860 -18626 -10826 -18586
rect -10786 -18626 -10770 -18586
rect -10930 -18660 -10770 -18626
rect -10930 -18700 -10900 -18660
rect -10860 -18700 -10826 -18660
rect -10786 -18700 -10770 -18660
rect -10930 -18730 -10770 -18700
rect -8930 -18586 -8770 -18560
rect -8930 -18626 -8900 -18586
rect -8860 -18626 -8826 -18586
rect -8786 -18626 -8770 -18586
rect -8930 -18660 -8770 -18626
rect -8930 -18700 -8900 -18660
rect -8860 -18700 -8826 -18660
rect -8786 -18700 -8770 -18660
rect -8930 -18730 -8770 -18700
rect -6930 -18586 -6770 -18560
rect -6930 -18626 -6900 -18586
rect -6860 -18626 -6826 -18586
rect -6786 -18626 -6770 -18586
rect -6930 -18660 -6770 -18626
rect -6930 -18700 -6900 -18660
rect -6860 -18700 -6826 -18660
rect -6786 -18700 -6770 -18660
rect -6930 -18730 -6770 -18700
rect -4930 -18586 -4770 -18560
rect -4930 -18626 -4900 -18586
rect -4860 -18626 -4826 -18586
rect -4786 -18626 -4770 -18586
rect -4930 -18660 -4770 -18626
rect -4930 -18700 -4900 -18660
rect -4860 -18700 -4826 -18660
rect -4786 -18700 -4770 -18660
rect -4930 -18730 -4770 -18700
rect -2930 -18586 -2770 -18560
rect -2930 -18626 -2900 -18586
rect -2860 -18626 -2826 -18586
rect -2786 -18626 -2770 -18586
rect -2930 -18660 -2770 -18626
rect -2930 -18700 -2900 -18660
rect -2860 -18700 -2826 -18660
rect -2786 -18700 -2770 -18660
rect -2930 -18730 -2770 -18700
rect -930 -18586 -770 -18560
rect -930 -18626 -900 -18586
rect -860 -18626 -826 -18586
rect -786 -18626 -770 -18586
rect -930 -18660 -770 -18626
rect -930 -18700 -900 -18660
rect -860 -18700 -826 -18660
rect -786 -18700 -770 -18660
rect -930 -18730 -770 -18700
rect 1070 -18586 1230 -18560
rect 1070 -18626 1100 -18586
rect 1140 -18626 1174 -18586
rect 1214 -18626 1230 -18586
rect 1070 -18660 1230 -18626
rect 1070 -18700 1100 -18660
rect 1140 -18700 1174 -18660
rect 1214 -18700 1230 -18660
rect 1070 -18730 1230 -18700
rect 3070 -18586 3230 -18560
rect 3070 -18626 3100 -18586
rect 3140 -18626 3174 -18586
rect 3214 -18626 3230 -18586
rect 3070 -18660 3230 -18626
rect 3070 -18700 3100 -18660
rect 3140 -18700 3174 -18660
rect 3214 -18700 3230 -18660
rect 3070 -18730 3230 -18700
rect 5070 -18586 5230 -18560
rect 5070 -18626 5100 -18586
rect 5140 -18626 5174 -18586
rect 5214 -18626 5230 -18586
rect 5070 -18660 5230 -18626
rect 5070 -18700 5100 -18660
rect 5140 -18700 5174 -18660
rect 5214 -18700 5230 -18660
rect 5070 -18730 5230 -18700
rect 7070 -18586 7230 -18560
rect 7070 -18626 7100 -18586
rect 7140 -18626 7174 -18586
rect 7214 -18626 7230 -18586
rect 7070 -18660 7230 -18626
rect 7070 -18700 7100 -18660
rect 7140 -18700 7174 -18660
rect 7214 -18700 7230 -18660
rect 7070 -18730 7230 -18700
rect 9070 -18586 9230 -18560
rect 9070 -18626 9100 -18586
rect 9140 -18626 9174 -18586
rect 9214 -18626 9230 -18586
rect 9070 -18660 9230 -18626
rect 9070 -18700 9100 -18660
rect 9140 -18700 9174 -18660
rect 9214 -18700 9230 -18660
rect 9070 -18730 9230 -18700
rect 11070 -18586 11230 -18560
rect 11070 -18626 11100 -18586
rect 11140 -18626 11174 -18586
rect 11214 -18626 11230 -18586
rect 11070 -18660 11230 -18626
rect 11070 -18700 11100 -18660
rect 11140 -18700 11174 -18660
rect 11214 -18700 11230 -18660
rect 11070 -18730 11230 -18700
rect 13070 -18586 13230 -18560
rect 13070 -18626 13100 -18586
rect 13140 -18626 13174 -18586
rect 13214 -18626 13230 -18586
rect 13070 -18660 13230 -18626
rect 13070 -18700 13100 -18660
rect 13140 -18700 13174 -18660
rect 13214 -18700 13230 -18660
rect 13070 -18730 13230 -18700
rect 15070 -18586 15230 -18560
rect 15070 -18626 15100 -18586
rect 15140 -18626 15174 -18586
rect 15214 -18626 15230 -18586
rect 15070 -18660 15230 -18626
rect 15070 -18700 15100 -18660
rect 15140 -18700 15174 -18660
rect 15214 -18700 15230 -18660
rect 15070 -18730 15230 -18700
rect 17070 -18586 17230 -18560
rect 17070 -18626 17100 -18586
rect 17140 -18626 17174 -18586
rect 17214 -18626 17230 -18586
rect 17070 -18660 17230 -18626
rect 17070 -18700 17100 -18660
rect 17140 -18700 17174 -18660
rect 17214 -18700 17230 -18660
rect 17070 -18730 17230 -18700
<< nsubdiffcont >>
rect -29880 24808 -29840 24848
rect -29806 24808 -29766 24848
rect -29880 24734 -29840 24774
rect -29806 24734 -29766 24774
rect -27880 24808 -27840 24848
rect -27806 24808 -27766 24848
rect -27880 24734 -27840 24774
rect -27806 24734 -27766 24774
rect -25880 24808 -25840 24848
rect -25806 24808 -25766 24848
rect -25880 24734 -25840 24774
rect -25806 24734 -25766 24774
rect -23880 24808 -23840 24848
rect -23806 24808 -23766 24848
rect -23880 24734 -23840 24774
rect -23806 24734 -23766 24774
rect -21880 24808 -21840 24848
rect -21806 24808 -21766 24848
rect -21880 24734 -21840 24774
rect -21806 24734 -21766 24774
rect -19880 24808 -19840 24848
rect -19806 24808 -19766 24848
rect -19880 24734 -19840 24774
rect -19806 24734 -19766 24774
rect -17880 24808 -17840 24848
rect -17806 24808 -17766 24848
rect -17880 24734 -17840 24774
rect -17806 24734 -17766 24774
rect -15880 24808 -15840 24848
rect -15806 24808 -15766 24848
rect -15880 24734 -15840 24774
rect -15806 24734 -15766 24774
rect -13880 24808 -13840 24848
rect -13806 24808 -13766 24848
rect -13880 24734 -13840 24774
rect -13806 24734 -13766 24774
rect -11880 24808 -11840 24848
rect -11806 24808 -11766 24848
rect -11880 24734 -11840 24774
rect -11806 24734 -11766 24774
rect -9880 24808 -9840 24848
rect -9806 24808 -9766 24848
rect -9880 24734 -9840 24774
rect -9806 24734 -9766 24774
rect -7880 24808 -7840 24848
rect -7806 24808 -7766 24848
rect -7880 24734 -7840 24774
rect -7806 24734 -7766 24774
rect -5880 24808 -5840 24848
rect -5806 24808 -5766 24848
rect -5880 24734 -5840 24774
rect -5806 24734 -5766 24774
rect -3880 24808 -3840 24848
rect -3806 24808 -3766 24848
rect -3880 24734 -3840 24774
rect -3806 24734 -3766 24774
rect -1880 24808 -1840 24848
rect -1806 24808 -1766 24848
rect -1880 24734 -1840 24774
rect -1806 24734 -1766 24774
rect 120 24808 160 24848
rect 194 24808 234 24848
rect 120 24734 160 24774
rect 194 24734 234 24774
rect 2120 24808 2160 24848
rect 2194 24808 2234 24848
rect 2120 24734 2160 24774
rect 2194 24734 2234 24774
rect 4120 24808 4160 24848
rect 4194 24808 4234 24848
rect 4120 24734 4160 24774
rect 4194 24734 4234 24774
rect 6120 24808 6160 24848
rect 6194 24808 6234 24848
rect 6120 24734 6160 24774
rect 6194 24734 6234 24774
rect 8120 24808 8160 24848
rect 8194 24808 8234 24848
rect 8120 24734 8160 24774
rect 8194 24734 8234 24774
rect 10120 24808 10160 24848
rect 10194 24808 10234 24848
rect 10120 24734 10160 24774
rect 10194 24734 10234 24774
rect 12120 24808 12160 24848
rect 12194 24808 12234 24848
rect 12120 24734 12160 24774
rect 12194 24734 12234 24774
rect 14120 24808 14160 24848
rect 14194 24808 14234 24848
rect 14120 24734 14160 24774
rect 14194 24734 14234 24774
rect 16120 24808 16160 24848
rect 16194 24808 16234 24848
rect 16120 24734 16160 24774
rect 16194 24734 16234 24774
rect 18120 24808 18160 24848
rect 18194 24808 18234 24848
rect 18120 24734 18160 24774
rect 18194 24734 18234 24774
rect 18250 24080 18290 24120
rect 18324 24080 18364 24120
rect 18250 24006 18290 24046
rect 18324 24006 18364 24046
rect -30086 23590 -30046 23630
rect -30012 23590 -29972 23630
rect -30086 23516 -30046 23556
rect -30012 23516 -29972 23556
rect 18250 22080 18290 22120
rect 18324 22080 18364 22120
rect 18250 22006 18290 22046
rect 18324 22006 18364 22046
rect -30086 21590 -30046 21630
rect -30012 21590 -29972 21630
rect -30086 21516 -30046 21556
rect -30012 21516 -29972 21556
rect 18250 20080 18290 20120
rect 18324 20080 18364 20120
rect 18250 20006 18290 20046
rect 18324 20006 18364 20046
rect -30086 19590 -30046 19630
rect -30012 19590 -29972 19630
rect -30086 19516 -30046 19556
rect -30012 19516 -29972 19556
rect 18250 18080 18290 18120
rect 18324 18080 18364 18120
rect 18250 18006 18290 18046
rect 18324 18006 18364 18046
rect -30086 17590 -30046 17630
rect -30012 17590 -29972 17630
rect -30086 17516 -30046 17556
rect -30012 17516 -29972 17556
rect 18250 16080 18290 16120
rect 18324 16080 18364 16120
rect 18250 16006 18290 16046
rect 18324 16006 18364 16046
rect -30086 15590 -30046 15630
rect -30012 15590 -29972 15630
rect -30086 15516 -30046 15556
rect -30012 15516 -29972 15556
rect 18250 14080 18290 14120
rect 18324 14080 18364 14120
rect 18250 14006 18290 14046
rect 18324 14006 18364 14046
rect -30086 13590 -30046 13630
rect -30012 13590 -29972 13630
rect -30086 13516 -30046 13556
rect -30012 13516 -29972 13556
rect 18250 12080 18290 12120
rect 18324 12080 18364 12120
rect 18250 12006 18290 12046
rect 18324 12006 18364 12046
rect -30086 11590 -30046 11630
rect -30012 11590 -29972 11630
rect -30086 11516 -30046 11556
rect -30012 11516 -29972 11556
rect 18250 10080 18290 10120
rect 18324 10080 18364 10120
rect 18250 10006 18290 10046
rect 18324 10006 18364 10046
rect -30086 9590 -30046 9630
rect -30012 9590 -29972 9630
rect -30086 9516 -30046 9556
rect -30012 9516 -29972 9556
rect 18250 8080 18290 8120
rect 18324 8080 18364 8120
rect 18250 8006 18290 8046
rect 18324 8006 18364 8046
rect -30086 7590 -30046 7630
rect -30012 7590 -29972 7630
rect -30086 7516 -30046 7556
rect -30012 7516 -29972 7556
rect 18250 6080 18290 6120
rect 18324 6080 18364 6120
rect 18250 6006 18290 6046
rect 18324 6006 18364 6046
rect -30086 5590 -30046 5630
rect -30012 5590 -29972 5630
rect -30086 5516 -30046 5556
rect -30012 5516 -29972 5556
rect 18250 4080 18290 4120
rect 18324 4080 18364 4120
rect 18250 4006 18290 4046
rect 18324 4006 18364 4046
rect -30086 3590 -30046 3630
rect -30012 3590 -29972 3630
rect -30086 3516 -30046 3556
rect -30012 3516 -29972 3556
rect 18250 2080 18290 2120
rect 18324 2080 18364 2120
rect 18250 2006 18290 2046
rect 18324 2006 18364 2046
rect -30086 1590 -30046 1630
rect -30012 1590 -29972 1630
rect -30086 1516 -30046 1556
rect -30012 1516 -29972 1556
rect 18250 80 18290 120
rect 18324 80 18364 120
rect 18250 6 18290 46
rect 18324 6 18364 46
rect -30086 -410 -30046 -370
rect -30012 -410 -29972 -370
rect -30086 -484 -30046 -444
rect -30012 -484 -29972 -444
rect 18250 -1920 18290 -1880
rect 18324 -1920 18364 -1880
rect 18250 -1994 18290 -1954
rect 18324 -1994 18364 -1954
rect -30086 -2410 -30046 -2370
rect -30012 -2410 -29972 -2370
rect -30086 -2484 -30046 -2444
rect -30012 -2484 -29972 -2444
rect 18250 -3920 18290 -3880
rect 18324 -3920 18364 -3880
rect 18250 -3994 18290 -3954
rect 18324 -3994 18364 -3954
rect -30086 -4410 -30046 -4370
rect -30012 -4410 -29972 -4370
rect -30086 -4484 -30046 -4444
rect -30012 -4484 -29972 -4444
rect 18250 -5920 18290 -5880
rect 18324 -5920 18364 -5880
rect 18250 -5994 18290 -5954
rect 18324 -5994 18364 -5954
rect -30086 -6410 -30046 -6370
rect -30012 -6410 -29972 -6370
rect -30086 -6484 -30046 -6444
rect -30012 -6484 -29972 -6444
rect 18250 -7920 18290 -7880
rect 18324 -7920 18364 -7880
rect 18250 -7994 18290 -7954
rect 18324 -7994 18364 -7954
rect -30086 -8410 -30046 -8370
rect -30012 -8410 -29972 -8370
rect -30086 -8484 -30046 -8444
rect -30012 -8484 -29972 -8444
rect 18250 -9920 18290 -9880
rect 18324 -9920 18364 -9880
rect 18250 -9994 18290 -9954
rect 18324 -9994 18364 -9954
rect -30086 -10410 -30046 -10370
rect -30012 -10410 -29972 -10370
rect -30086 -10484 -30046 -10444
rect -30012 -10484 -29972 -10444
rect 18250 -11920 18290 -11880
rect 18324 -11920 18364 -11880
rect 18250 -11994 18290 -11954
rect 18324 -11994 18364 -11954
rect -30086 -12410 -30046 -12370
rect -30012 -12410 -29972 -12370
rect -30086 -12484 -30046 -12444
rect -30012 -12484 -29972 -12444
rect 18250 -13920 18290 -13880
rect 18324 -13920 18364 -13880
rect 18250 -13994 18290 -13954
rect 18324 -13994 18364 -13954
rect -30086 -14410 -30046 -14370
rect -30012 -14410 -29972 -14370
rect -30086 -14484 -30046 -14444
rect -30012 -14484 -29972 -14444
rect 18250 -15920 18290 -15880
rect 18324 -15920 18364 -15880
rect 18250 -15994 18290 -15954
rect 18324 -15994 18364 -15954
rect -30086 -16410 -30046 -16370
rect -30012 -16410 -29972 -16370
rect -30086 -16484 -30046 -16444
rect -30012 -16484 -29972 -16444
rect 18250 -17920 18290 -17880
rect 18324 -17920 18364 -17880
rect 18250 -17994 18290 -17954
rect 18324 -17994 18364 -17954
rect -30086 -18410 -30046 -18370
rect -30012 -18410 -29972 -18370
rect -30086 -18484 -30046 -18444
rect -30012 -18484 -29972 -18444
rect -28900 -18626 -28860 -18586
rect -28826 -18626 -28786 -18586
rect -28900 -18700 -28860 -18660
rect -28826 -18700 -28786 -18660
rect -26900 -18626 -26860 -18586
rect -26826 -18626 -26786 -18586
rect -26900 -18700 -26860 -18660
rect -26826 -18700 -26786 -18660
rect -24900 -18626 -24860 -18586
rect -24826 -18626 -24786 -18586
rect -24900 -18700 -24860 -18660
rect -24826 -18700 -24786 -18660
rect -22900 -18626 -22860 -18586
rect -22826 -18626 -22786 -18586
rect -22900 -18700 -22860 -18660
rect -22826 -18700 -22786 -18660
rect -20900 -18626 -20860 -18586
rect -20826 -18626 -20786 -18586
rect -20900 -18700 -20860 -18660
rect -20826 -18700 -20786 -18660
rect -18900 -18626 -18860 -18586
rect -18826 -18626 -18786 -18586
rect -18900 -18700 -18860 -18660
rect -18826 -18700 -18786 -18660
rect -16900 -18626 -16860 -18586
rect -16826 -18626 -16786 -18586
rect -16900 -18700 -16860 -18660
rect -16826 -18700 -16786 -18660
rect -14900 -18626 -14860 -18586
rect -14826 -18626 -14786 -18586
rect -14900 -18700 -14860 -18660
rect -14826 -18700 -14786 -18660
rect -12900 -18626 -12860 -18586
rect -12826 -18626 -12786 -18586
rect -12900 -18700 -12860 -18660
rect -12826 -18700 -12786 -18660
rect -10900 -18626 -10860 -18586
rect -10826 -18626 -10786 -18586
rect -10900 -18700 -10860 -18660
rect -10826 -18700 -10786 -18660
rect -8900 -18626 -8860 -18586
rect -8826 -18626 -8786 -18586
rect -8900 -18700 -8860 -18660
rect -8826 -18700 -8786 -18660
rect -6900 -18626 -6860 -18586
rect -6826 -18626 -6786 -18586
rect -6900 -18700 -6860 -18660
rect -6826 -18700 -6786 -18660
rect -4900 -18626 -4860 -18586
rect -4826 -18626 -4786 -18586
rect -4900 -18700 -4860 -18660
rect -4826 -18700 -4786 -18660
rect -2900 -18626 -2860 -18586
rect -2826 -18626 -2786 -18586
rect -2900 -18700 -2860 -18660
rect -2826 -18700 -2786 -18660
rect -900 -18626 -860 -18586
rect -826 -18626 -786 -18586
rect -900 -18700 -860 -18660
rect -826 -18700 -786 -18660
rect 1100 -18626 1140 -18586
rect 1174 -18626 1214 -18586
rect 1100 -18700 1140 -18660
rect 1174 -18700 1214 -18660
rect 3100 -18626 3140 -18586
rect 3174 -18626 3214 -18586
rect 3100 -18700 3140 -18660
rect 3174 -18700 3214 -18660
rect 5100 -18626 5140 -18586
rect 5174 -18626 5214 -18586
rect 5100 -18700 5140 -18660
rect 5174 -18700 5214 -18660
rect 7100 -18626 7140 -18586
rect 7174 -18626 7214 -18586
rect 7100 -18700 7140 -18660
rect 7174 -18700 7214 -18660
rect 9100 -18626 9140 -18586
rect 9174 -18626 9214 -18586
rect 9100 -18700 9140 -18660
rect 9174 -18700 9214 -18660
rect 11100 -18626 11140 -18586
rect 11174 -18626 11214 -18586
rect 11100 -18700 11140 -18660
rect 11174 -18700 11214 -18660
rect 13100 -18626 13140 -18586
rect 13174 -18626 13214 -18586
rect 13100 -18700 13140 -18660
rect 13174 -18700 13214 -18660
rect 15100 -18626 15140 -18586
rect 15174 -18626 15214 -18586
rect 15100 -18700 15140 -18660
rect 15174 -18700 15214 -18660
rect 17100 -18626 17140 -18586
rect 17174 -18626 17214 -18586
rect 17100 -18700 17140 -18660
rect 17174 -18700 17214 -18660
<< locali >>
rect -30116 24848 18381 24874
rect -30116 24808 -29880 24848
rect -29840 24808 -29806 24848
rect -29766 24808 -27880 24848
rect -27840 24808 -27806 24848
rect -27766 24808 -25880 24848
rect -25840 24808 -25806 24848
rect -25766 24808 -23880 24848
rect -23840 24808 -23806 24848
rect -23766 24808 -21880 24848
rect -21840 24808 -21806 24848
rect -21766 24808 -19880 24848
rect -19840 24808 -19806 24848
rect -19766 24808 -17880 24848
rect -17840 24808 -17806 24848
rect -17766 24808 -15880 24848
rect -15840 24808 -15806 24848
rect -15766 24808 -13880 24848
rect -13840 24808 -13806 24848
rect -13766 24808 -11880 24848
rect -11840 24808 -11806 24848
rect -11766 24808 -9880 24848
rect -9840 24808 -9806 24848
rect -9766 24808 -7880 24848
rect -7840 24808 -7806 24848
rect -7766 24808 -5880 24848
rect -5840 24808 -5806 24848
rect -5766 24808 -3880 24848
rect -3840 24808 -3806 24848
rect -3766 24808 -1880 24848
rect -1840 24808 -1806 24848
rect -1766 24808 120 24848
rect 160 24808 194 24848
rect 234 24808 2120 24848
rect 2160 24808 2194 24848
rect 2234 24808 4120 24848
rect 4160 24808 4194 24848
rect 4234 24808 6120 24848
rect 6160 24808 6194 24848
rect 6234 24808 8120 24848
rect 8160 24808 8194 24848
rect 8234 24808 10120 24848
rect 10160 24808 10194 24848
rect 10234 24808 12120 24848
rect 12160 24808 12194 24848
rect 12234 24808 14120 24848
rect 14160 24808 14194 24848
rect 14234 24808 16120 24848
rect 16160 24808 16194 24848
rect 16234 24808 18120 24848
rect 18160 24808 18194 24848
rect 18234 24808 18381 24848
rect -30116 24774 18381 24808
rect -30116 24734 -29880 24774
rect -29840 24734 -29806 24774
rect -29766 24734 -27880 24774
rect -27840 24734 -27806 24774
rect -27766 24734 -25880 24774
rect -25840 24734 -25806 24774
rect -25766 24734 -23880 24774
rect -23840 24734 -23806 24774
rect -23766 24734 -21880 24774
rect -21840 24734 -21806 24774
rect -21766 24734 -19880 24774
rect -19840 24734 -19806 24774
rect -19766 24734 -17880 24774
rect -17840 24734 -17806 24774
rect -17766 24734 -15880 24774
rect -15840 24734 -15806 24774
rect -15766 24734 -13880 24774
rect -13840 24734 -13806 24774
rect -13766 24734 -11880 24774
rect -11840 24734 -11806 24774
rect -11766 24734 -9880 24774
rect -9840 24734 -9806 24774
rect -9766 24734 -7880 24774
rect -7840 24734 -7806 24774
rect -7766 24734 -5880 24774
rect -5840 24734 -5806 24774
rect -5766 24734 -3880 24774
rect -3840 24734 -3806 24774
rect -3766 24734 -1880 24774
rect -1840 24734 -1806 24774
rect -1766 24734 120 24774
rect 160 24734 194 24774
rect 234 24734 2120 24774
rect 2160 24734 2194 24774
rect 2234 24734 4120 24774
rect 4160 24734 4194 24774
rect 4234 24734 6120 24774
rect 6160 24734 6194 24774
rect 6234 24734 8120 24774
rect 8160 24734 8194 24774
rect 8234 24734 10120 24774
rect 10160 24734 10194 24774
rect 10234 24734 12120 24774
rect 12160 24734 12194 24774
rect 12234 24734 14120 24774
rect 14160 24734 14194 24774
rect 14234 24734 16120 24774
rect 16160 24734 16194 24774
rect 16234 24734 18120 24774
rect 18160 24734 18194 24774
rect 18234 24734 18381 24774
rect -30116 24668 18381 24734
rect -30116 23630 -29910 24668
rect -30116 23590 -30086 23630
rect -30046 23590 -30012 23630
rect -29972 23590 -29910 23630
rect -30116 23556 -29910 23590
rect -30116 23516 -30086 23556
rect -30046 23516 -30012 23556
rect -29972 23516 -29910 23556
rect -30116 21630 -29910 23516
rect -30116 21590 -30086 21630
rect -30046 21590 -30012 21630
rect -29972 21590 -29910 21630
rect -30116 21556 -29910 21590
rect -30116 21516 -30086 21556
rect -30046 21516 -30012 21556
rect -29972 21516 -29910 21556
rect -30116 19630 -29910 21516
rect -30116 19590 -30086 19630
rect -30046 19590 -30012 19630
rect -29972 19590 -29910 19630
rect -30116 19556 -29910 19590
rect -30116 19516 -30086 19556
rect -30046 19516 -30012 19556
rect -29972 19516 -29910 19556
rect -30116 17630 -29910 19516
rect -30116 17590 -30086 17630
rect -30046 17590 -30012 17630
rect -29972 17590 -29910 17630
rect -30116 17556 -29910 17590
rect -30116 17516 -30086 17556
rect -30046 17516 -30012 17556
rect -29972 17516 -29910 17556
rect -30116 15630 -29910 17516
rect -30116 15590 -30086 15630
rect -30046 15590 -30012 15630
rect -29972 15590 -29910 15630
rect -30116 15556 -29910 15590
rect -30116 15516 -30086 15556
rect -30046 15516 -30012 15556
rect -29972 15516 -29910 15556
rect -30116 13630 -29910 15516
rect -30116 13590 -30086 13630
rect -30046 13590 -30012 13630
rect -29972 13590 -29910 13630
rect -30116 13556 -29910 13590
rect -30116 13516 -30086 13556
rect -30046 13516 -30012 13556
rect -29972 13516 -29910 13556
rect -30116 11630 -29910 13516
rect -30116 11590 -30086 11630
rect -30046 11590 -30012 11630
rect -29972 11590 -29910 11630
rect -30116 11556 -29910 11590
rect -30116 11516 -30086 11556
rect -30046 11516 -30012 11556
rect -29972 11516 -29910 11556
rect -30116 9630 -29910 11516
rect -30116 9590 -30086 9630
rect -30046 9590 -30012 9630
rect -29972 9590 -29910 9630
rect -30116 9556 -29910 9590
rect -30116 9516 -30086 9556
rect -30046 9516 -30012 9556
rect -29972 9516 -29910 9556
rect -30116 7630 -29910 9516
rect -30116 7590 -30086 7630
rect -30046 7590 -30012 7630
rect -29972 7590 -29910 7630
rect -30116 7556 -29910 7590
rect -30116 7516 -30086 7556
rect -30046 7516 -30012 7556
rect -29972 7516 -29910 7556
rect -30116 5630 -29910 7516
rect -30116 5590 -30086 5630
rect -30046 5590 -30012 5630
rect -29972 5590 -29910 5630
rect -30116 5556 -29910 5590
rect -30116 5516 -30086 5556
rect -30046 5516 -30012 5556
rect -29972 5516 -29910 5556
rect -30116 3630 -29910 5516
rect -30116 3590 -30086 3630
rect -30046 3590 -30012 3630
rect -29972 3590 -29910 3630
rect -30116 3556 -29910 3590
rect -30116 3516 -30086 3556
rect -30046 3516 -30012 3556
rect -29972 3516 -29910 3556
rect -30116 1630 -29910 3516
rect -30116 1590 -30086 1630
rect -30046 1590 -30012 1630
rect -29972 1590 -29910 1630
rect -30116 1556 -29910 1590
rect -30116 1516 -30086 1556
rect -30046 1516 -30012 1556
rect -29972 1516 -29910 1556
rect -30116 -370 -29910 1516
rect -30116 -410 -30086 -370
rect -30046 -410 -30012 -370
rect -29972 -410 -29910 -370
rect -30116 -444 -29910 -410
rect -30116 -484 -30086 -444
rect -30046 -484 -30012 -444
rect -29972 -484 -29910 -444
rect -30116 -2370 -29910 -484
rect -30116 -2410 -30086 -2370
rect -30046 -2410 -30012 -2370
rect -29972 -2410 -29910 -2370
rect -30116 -2444 -29910 -2410
rect -30116 -2484 -30086 -2444
rect -30046 -2484 -30012 -2444
rect -29972 -2484 -29910 -2444
rect -30116 -4370 -29910 -2484
rect -30116 -4410 -30086 -4370
rect -30046 -4410 -30012 -4370
rect -29972 -4410 -29910 -4370
rect -30116 -4444 -29910 -4410
rect -30116 -4484 -30086 -4444
rect -30046 -4484 -30012 -4444
rect -29972 -4484 -29910 -4444
rect -30116 -6370 -29910 -4484
rect -30116 -6410 -30086 -6370
rect -30046 -6410 -30012 -6370
rect -29972 -6410 -29910 -6370
rect -30116 -6444 -29910 -6410
rect -30116 -6484 -30086 -6444
rect -30046 -6484 -30012 -6444
rect -29972 -6484 -29910 -6444
rect -30116 -8370 -29910 -6484
rect -30116 -8410 -30086 -8370
rect -30046 -8410 -30012 -8370
rect -29972 -8410 -29910 -8370
rect -30116 -8444 -29910 -8410
rect -30116 -8484 -30086 -8444
rect -30046 -8484 -30012 -8444
rect -29972 -8484 -29910 -8444
rect -30116 -10370 -29910 -8484
rect -30116 -10410 -30086 -10370
rect -30046 -10410 -30012 -10370
rect -29972 -10410 -29910 -10370
rect -30116 -10444 -29910 -10410
rect -30116 -10484 -30086 -10444
rect -30046 -10484 -30012 -10444
rect -29972 -10484 -29910 -10444
rect -30116 -12370 -29910 -10484
rect -30116 -12410 -30086 -12370
rect -30046 -12410 -30012 -12370
rect -29972 -12410 -29910 -12370
rect -30116 -12444 -29910 -12410
rect -30116 -12484 -30086 -12444
rect -30046 -12484 -30012 -12444
rect -29972 -12484 -29910 -12444
rect -30116 -14370 -29910 -12484
rect -30116 -14410 -30086 -14370
rect -30046 -14410 -30012 -14370
rect -29972 -14410 -29910 -14370
rect -30116 -14444 -29910 -14410
rect -30116 -14484 -30086 -14444
rect -30046 -14484 -30012 -14444
rect -29972 -14484 -29910 -14444
rect -30116 -16370 -29910 -14484
rect -30116 -16410 -30086 -16370
rect -30046 -16410 -30012 -16370
rect -29972 -16410 -29910 -16370
rect -30116 -16444 -29910 -16410
rect -30116 -16484 -30086 -16444
rect -30046 -16484 -30012 -16444
rect -29972 -16484 -29910 -16444
rect -30116 -18370 -29910 -16484
rect -30116 -18410 -30086 -18370
rect -30046 -18410 -30012 -18370
rect -29972 -18410 -29910 -18370
rect -30116 -18444 -29910 -18410
rect -30116 -18484 -30086 -18444
rect -30046 -18484 -30012 -18444
rect -29972 -18484 -29910 -18444
rect -30116 -18524 -29910 -18484
rect 18175 24120 18381 24668
rect 18175 24080 18250 24120
rect 18290 24080 18324 24120
rect 18364 24080 18381 24120
rect 18175 24046 18381 24080
rect 18175 24006 18250 24046
rect 18290 24006 18324 24046
rect 18364 24006 18381 24046
rect 18175 22120 18381 24006
rect 18175 22080 18250 22120
rect 18290 22080 18324 22120
rect 18364 22080 18381 22120
rect 18175 22046 18381 22080
rect 18175 22006 18250 22046
rect 18290 22006 18324 22046
rect 18364 22006 18381 22046
rect 18175 20120 18381 22006
rect 18175 20080 18250 20120
rect 18290 20080 18324 20120
rect 18364 20080 18381 20120
rect 18175 20046 18381 20080
rect 18175 20006 18250 20046
rect 18290 20006 18324 20046
rect 18364 20006 18381 20046
rect 18175 18120 18381 20006
rect 18175 18080 18250 18120
rect 18290 18080 18324 18120
rect 18364 18080 18381 18120
rect 18175 18046 18381 18080
rect 18175 18006 18250 18046
rect 18290 18006 18324 18046
rect 18364 18006 18381 18046
rect 18175 16120 18381 18006
rect 18175 16080 18250 16120
rect 18290 16080 18324 16120
rect 18364 16080 18381 16120
rect 18175 16046 18381 16080
rect 18175 16006 18250 16046
rect 18290 16006 18324 16046
rect 18364 16006 18381 16046
rect 18175 14120 18381 16006
rect 18175 14080 18250 14120
rect 18290 14080 18324 14120
rect 18364 14080 18381 14120
rect 18175 14046 18381 14080
rect 18175 14006 18250 14046
rect 18290 14006 18324 14046
rect 18364 14006 18381 14046
rect 18175 12120 18381 14006
rect 18175 12080 18250 12120
rect 18290 12080 18324 12120
rect 18364 12080 18381 12120
rect 18175 12046 18381 12080
rect 18175 12006 18250 12046
rect 18290 12006 18324 12046
rect 18364 12006 18381 12046
rect 18175 10120 18381 12006
rect 18175 10080 18250 10120
rect 18290 10080 18324 10120
rect 18364 10080 18381 10120
rect 18175 10046 18381 10080
rect 18175 10006 18250 10046
rect 18290 10006 18324 10046
rect 18364 10006 18381 10046
rect 18175 8120 18381 10006
rect 18175 8080 18250 8120
rect 18290 8080 18324 8120
rect 18364 8080 18381 8120
rect 18175 8046 18381 8080
rect 18175 8006 18250 8046
rect 18290 8006 18324 8046
rect 18364 8006 18381 8046
rect 18175 6120 18381 8006
rect 18175 6080 18250 6120
rect 18290 6080 18324 6120
rect 18364 6080 18381 6120
rect 18175 6046 18381 6080
rect 18175 6006 18250 6046
rect 18290 6006 18324 6046
rect 18364 6006 18381 6046
rect 18175 4120 18381 6006
rect 18175 4080 18250 4120
rect 18290 4080 18324 4120
rect 18364 4080 18381 4120
rect 18175 4046 18381 4080
rect 18175 4006 18250 4046
rect 18290 4006 18324 4046
rect 18364 4006 18381 4046
rect 18175 2120 18381 4006
rect 18175 2080 18250 2120
rect 18290 2080 18324 2120
rect 18364 2080 18381 2120
rect 18175 2046 18381 2080
rect 18175 2006 18250 2046
rect 18290 2006 18324 2046
rect 18364 2006 18381 2046
rect 18175 120 18381 2006
rect 18175 80 18250 120
rect 18290 80 18324 120
rect 18364 80 18381 120
rect 18175 46 18381 80
rect 18175 6 18250 46
rect 18290 6 18324 46
rect 18364 6 18381 46
rect 18175 -1880 18381 6
rect 18175 -1920 18250 -1880
rect 18290 -1920 18324 -1880
rect 18364 -1920 18381 -1880
rect 18175 -1954 18381 -1920
rect 18175 -1994 18250 -1954
rect 18290 -1994 18324 -1954
rect 18364 -1994 18381 -1954
rect 18175 -3880 18381 -1994
rect 18175 -3920 18250 -3880
rect 18290 -3920 18324 -3880
rect 18364 -3920 18381 -3880
rect 18175 -3954 18381 -3920
rect 18175 -3994 18250 -3954
rect 18290 -3994 18324 -3954
rect 18364 -3994 18381 -3954
rect 18175 -5880 18381 -3994
rect 18175 -5920 18250 -5880
rect 18290 -5920 18324 -5880
rect 18364 -5920 18381 -5880
rect 18175 -5954 18381 -5920
rect 18175 -5994 18250 -5954
rect 18290 -5994 18324 -5954
rect 18364 -5994 18381 -5954
rect 18175 -7880 18381 -5994
rect 18175 -7920 18250 -7880
rect 18290 -7920 18324 -7880
rect 18364 -7920 18381 -7880
rect 18175 -7954 18381 -7920
rect 18175 -7994 18250 -7954
rect 18290 -7994 18324 -7954
rect 18364 -7994 18381 -7954
rect 18175 -9880 18381 -7994
rect 18175 -9920 18250 -9880
rect 18290 -9920 18324 -9880
rect 18364 -9920 18381 -9880
rect 18175 -9954 18381 -9920
rect 18175 -9994 18250 -9954
rect 18290 -9994 18324 -9954
rect 18364 -9994 18381 -9954
rect 18175 -11880 18381 -9994
rect 18175 -11920 18250 -11880
rect 18290 -11920 18324 -11880
rect 18364 -11920 18381 -11880
rect 18175 -11954 18381 -11920
rect 18175 -11994 18250 -11954
rect 18290 -11994 18324 -11954
rect 18364 -11994 18381 -11954
rect 18175 -13880 18381 -11994
rect 18175 -13920 18250 -13880
rect 18290 -13920 18324 -13880
rect 18364 -13920 18381 -13880
rect 18175 -13954 18381 -13920
rect 18175 -13994 18250 -13954
rect 18290 -13994 18324 -13954
rect 18364 -13994 18381 -13954
rect 18175 -15880 18381 -13994
rect 18175 -15920 18250 -15880
rect 18290 -15920 18324 -15880
rect 18364 -15920 18381 -15880
rect 18175 -15954 18381 -15920
rect 18175 -15994 18250 -15954
rect 18290 -15994 18324 -15954
rect 18364 -15994 18381 -15954
rect 18175 -17880 18381 -15994
rect 18175 -17920 18250 -17880
rect 18290 -17920 18324 -17880
rect 18364 -17920 18381 -17880
rect 18175 -17954 18381 -17920
rect 18175 -17994 18250 -17954
rect 18290 -17994 18324 -17954
rect 18364 -17994 18381 -17954
rect 18175 -18524 18381 -17994
rect -30116 -18586 18381 -18524
rect -30116 -18626 -28900 -18586
rect -28860 -18626 -28826 -18586
rect -28786 -18626 -26900 -18586
rect -26860 -18626 -26826 -18586
rect -26786 -18626 -24900 -18586
rect -24860 -18626 -24826 -18586
rect -24786 -18626 -22900 -18586
rect -22860 -18626 -22826 -18586
rect -22786 -18626 -20900 -18586
rect -20860 -18626 -20826 -18586
rect -20786 -18626 -18900 -18586
rect -18860 -18626 -18826 -18586
rect -18786 -18626 -16900 -18586
rect -16860 -18626 -16826 -18586
rect -16786 -18626 -14900 -18586
rect -14860 -18626 -14826 -18586
rect -14786 -18626 -12900 -18586
rect -12860 -18626 -12826 -18586
rect -12786 -18626 -10900 -18586
rect -10860 -18626 -10826 -18586
rect -10786 -18626 -8900 -18586
rect -8860 -18626 -8826 -18586
rect -8786 -18626 -6900 -18586
rect -6860 -18626 -6826 -18586
rect -6786 -18626 -4900 -18586
rect -4860 -18626 -4826 -18586
rect -4786 -18626 -2900 -18586
rect -2860 -18626 -2826 -18586
rect -2786 -18626 -900 -18586
rect -860 -18626 -826 -18586
rect -786 -18626 1100 -18586
rect 1140 -18626 1174 -18586
rect 1214 -18626 3100 -18586
rect 3140 -18626 3174 -18586
rect 3214 -18626 5100 -18586
rect 5140 -18626 5174 -18586
rect 5214 -18626 7100 -18586
rect 7140 -18626 7174 -18586
rect 7214 -18626 9100 -18586
rect 9140 -18626 9174 -18586
rect 9214 -18626 11100 -18586
rect 11140 -18626 11174 -18586
rect 11214 -18626 13100 -18586
rect 13140 -18626 13174 -18586
rect 13214 -18626 15100 -18586
rect 15140 -18626 15174 -18586
rect 15214 -18626 17100 -18586
rect 17140 -18626 17174 -18586
rect 17214 -18626 18381 -18586
rect -30116 -18660 18381 -18626
rect -30116 -18700 -28900 -18660
rect -28860 -18700 -28826 -18660
rect -28786 -18700 -26900 -18660
rect -26860 -18700 -26826 -18660
rect -26786 -18700 -24900 -18660
rect -24860 -18700 -24826 -18660
rect -24786 -18700 -22900 -18660
rect -22860 -18700 -22826 -18660
rect -22786 -18700 -20900 -18660
rect -20860 -18700 -20826 -18660
rect -20786 -18700 -18900 -18660
rect -18860 -18700 -18826 -18660
rect -18786 -18700 -16900 -18660
rect -16860 -18700 -16826 -18660
rect -16786 -18700 -14900 -18660
rect -14860 -18700 -14826 -18660
rect -14786 -18700 -12900 -18660
rect -12860 -18700 -12826 -18660
rect -12786 -18700 -10900 -18660
rect -10860 -18700 -10826 -18660
rect -10786 -18700 -8900 -18660
rect -8860 -18700 -8826 -18660
rect -8786 -18700 -6900 -18660
rect -6860 -18700 -6826 -18660
rect -6786 -18700 -4900 -18660
rect -4860 -18700 -4826 -18660
rect -4786 -18700 -2900 -18660
rect -2860 -18700 -2826 -18660
rect -2786 -18700 -900 -18660
rect -860 -18700 -826 -18660
rect -786 -18700 1100 -18660
rect 1140 -18700 1174 -18660
rect 1214 -18700 3100 -18660
rect 3140 -18700 3174 -18660
rect 3214 -18700 5100 -18660
rect 5140 -18700 5174 -18660
rect 5214 -18700 7100 -18660
rect 7140 -18700 7174 -18660
rect 7214 -18700 9100 -18660
rect 9140 -18700 9174 -18660
rect 9214 -18700 11100 -18660
rect 11140 -18700 11174 -18660
rect 11214 -18700 13100 -18660
rect 13140 -18700 13174 -18660
rect 13214 -18700 15100 -18660
rect 15140 -18700 15174 -18660
rect 15214 -18700 17100 -18660
rect 17140 -18700 17174 -18660
rect 17214 -18700 18381 -18660
rect -30116 -18730 18381 -18700
<< metal1 >>
rect -30116 24668 18381 24874
rect -30116 -18524 -29910 24668
rect -3328 -16710 -2408 -16590
rect -3328 -18017 -3208 -16710
rect -9902 -18083 -3208 -18017
rect 18175 -18524 18381 24668
rect -30116 -18730 18381 -18524
<< metal2 >>
rect -11563 -7342 -11363 -4237
rect -11563 -7462 -2412 -7342
rect -3208 -16710 -2408 -16590
use ONES_COUNTER  ONES_COUNTER_0
timestamp 1713591521
transform 1 0 -3101 0 1 -18207
box 0 824 11908 12912
use SDC  SDC_0
timestamp 1713591521
transform 1 0 19 0 1 -21
box -29735 -18309 17962 24495
<< end >>
