* NGSPICE file created from ONES_COUNTER_pex.ext - technology: sky130A

.subckt ONES_COUNTER_pex VGND VPWR clk rst pulse ready ones[0] ones[1] ones[2] ones[3] ones[4] ones[5]
+ ones[6] ones[7] ones[8] ones[9] ones[10]
X0 _067_ a_5363_2880# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=135.43779 ps=1.28947k w=0.87 l=1.05
X2 VPWR a_2823_4943# a_2991_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X3 a_8999_5639# a_9095_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VGND a_7407_4667# a_7365_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X5 a_9213_3463# counter\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X6 VPWR a_3697_6031# a_3797_6147# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X7 a_6169_6549# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 a_2907_4943# a_2125_4949# a_2823_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_3053_8751# net6 a_2971_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X11 _049_ a_1670_6351# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 a_9163_3855# a_8381_3861# a_9079_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=87.036446 ps=919.38995 w=0.55 l=2.89
X14 net7 a_4279_2741# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 a_5837_5303# _059_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.122275 ps=1.08 w=0.42 l=0.15
X16 VPWR a_5142_3423# a_5069_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X17 VGND _068_ a_3273_2251# VGND sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VGND a_9919_4087# _033_ VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X19 VPWR a_8643_6249# a_8650_6153# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X20 a_4697_5461# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X21 VGND counter\[10\] a_5537_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X23 _039_ a_7663_7485# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X24 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X25 a_4709_5309# _060_ a_4627_5056# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X26 a_7290_7119# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X27 a_9677_3311# counter\[1\] _062_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X28 VGND a_2807_7093# a_2765_7497# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X29 a_4307_8439# a_4580_8439# a_4538_8567# VGND sky130_fd_pr__nfet_01v8 ad=0.107825 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 a_7369_9117# a_6835_8751# a_7274_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X31 a_8338_11177# _068_ a_8256_11177# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 a_2668_4405# _060_ a_2596_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X33 VGND net4 _052_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 a_5418_4511# a_5250_4765# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X35 a_6633_5487# a_6467_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X36 a_7791_9295# a_7093_9301# a_7534_9269# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X37 a_9832_8181# counter\[1\] a_10055_8527# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X38 a_9379_5461# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X39 VGND _025_ _012_ VGND sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
X40 a_10199_3285# pulse VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X41 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X42 VGND a_6169_6549# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X43 clknet_0_clk a_6169_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X44 VGND a_6423_11079# _057_ VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X45 a_9845_3087# net12 a_10039_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X46 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X47 VPWR clknet_1_0__leaf_clk a_3247_2773# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X48 VGND _093_ _011_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X49 a_10199_2197# rst VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X50 a_5801_4399# a_4811_4399# a_5675_4765# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X51 VPWR _068_ a_1499_5056# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X52 a_3697_6031# _080_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X53 VPWR a_4771_2741# _055_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X54 a_9586_5461# a_9386_5761# a_9735_5487# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X55 clknet_1_1__leaf_clk a_8390_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X56 a_6814_4765# a_6541_4399# a_6729_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X57 VGND _037_ a_7939_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X58 _081_ a_2682_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X59 VPWR a_4697_5461# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X60 _012_ _024_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.112125 ps=0.995 w=0.65 l=0.15
X61 a_7093_9301# a_6927_9301# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X62 VPWR a_4595_4073# a_4602_3977# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X63 _052_ net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X64 _030_ a_7980_4649# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X65 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X66 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X67 a_8381_3861# a_8215_3861# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X68 a_9586_5461# a_9379_5461# a_9762_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X69 a_9558_4917# a_9390_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X70 VGND a_9832_8181# _069_ VGND sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X71 a_9933_5487# a_9379_5461# a_9586_5461# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X72 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X73 a_9325_8573# _077_ a_9253_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X74 a_2398_4943# a_1959_4949# a_2313_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X75 a_9117_4949# a_8951_4949# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X76 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X77 a_6003_10089# counter\[2\] a_5785_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X78 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X79 a_9762_5853# a_9515_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X80 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X81 a_8215_10496# _030_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X82 VGND _010_ a_9197_6409# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X83 a_8601_6031# a_8263_6263# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X84 ones[3] a_10239_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X85 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X86 a_6475_7913# a_6283_7669# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X87 a_9961_8527# counter\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X88 a_2046_6575# a_1731_6727# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X89 VGND a_8390_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X90 VGND a_2639_7119# a_2807_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X91 a_3854_2741# a_3686_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X92 VPWR a_6982_4511# a_6909_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X93 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X94 counter\[2\] a_6719_10615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X95 a_6446_3677# a_6173_3311# a_6361_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X96 a_2524_5321# a_2125_4949# a_2398_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X97 a_4229_10761# a_3682_10505# a_3882_10660# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X98 a_2555_10704# counter\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X99 a_5169_3133# counter\[4\] a_5063_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X100 a_6515_4074# _029_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X101 a_2409_4445# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X102 VGND net2 a_9096_4373# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X103 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X104 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X105 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X106 VPWR _034_ a_2697_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X107 a_7074_5599# a_6906_5853# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X108 a_9896_9001# _084_ a_9435_9001# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
X109 a_3799_10927# _071_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X110 a_9314_5487# a_8999_5639# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X111 a_6541_6037# a_6375_6037# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X112 a_7074_5599# a_6906_5853# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X113 VGND a_4697_5461# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X114 VPWR _031_ a_6557_7913# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X115 a_4078_8757# _060_ a_3997_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.05355 ps=0.675 w=0.42 l=0.15
X116 a_6425_10602# _045_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X117 VPWR a_7791_9295# a_7959_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X119 a_6719_10615# a_6887_10615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X120 VGND a_8822_3829# a_8780_4233# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X121 a_9933_5487# a_9386_5761# a_9586_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X122 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X123 a_2125_4949# a_1959_4949# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X124 a_7366_9295# a_6927_9301# a_7281_9295# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X125 VPWR net9 a_10239_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X126 VPWR _046_ a_8447_5175# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X127 a_7171_10601# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X128 VGND clk a_6169_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X129 a_8390_7119# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X131 VGND a_4981_9991# _023_ VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X132 VPWR a_8631_2986# _014_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X133 a_7875_9295# a_7093_9301# a_7791_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X134 VPWR a_6614_3423# a_6541_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X135 VPWR clknet_0_clk a_4697_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X136 VGND counter\[6\] a_4668_7913# VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X137 clknet_1_0__leaf_clk a_4697_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X138 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X139 _088_ a_2460_3971# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X140 VPWR a_5843_4667# counter\[0\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X141 a_7492_9673# a_7093_9301# a_7366_9295# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X142 VPWR net1 a_7290_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X143 VGND net3 a_10239_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X144 _084_ counter\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X145 a_4311_4087# a_4595_4073# a_4530_4221# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X146 a_6541_3677# a_6007_3311# a_6446_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X147 VGND a_3854_2741# a_3812_3145# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X148 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X149 VPWR _054_ a_5087_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X150 a_7725_10761# a_7171_10601# a_7378_10660# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X151 a_6982_6005# a_6814_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X152 clknet_0_clk a_6169_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X153 VPWR a_6169_6549# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X154 a_8569_3855# _015_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X155 _050_ net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X156 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X157 a_3633_10383# a_3295_10615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X158 VPWR clknet_1_1__leaf_clk a_6927_9301# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X159 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X160 VPWR _028_ a_8215_10496# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X161 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X162 VGND a_8907_2986# _008_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X163 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X164 a_6703_2197# a_6987_2197# a_6922_2223# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X165 VGND net9 a_10239_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X166 net14 a_7867_9019# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X167 a_8113_2223# counter\[1\] _065_ VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X168 a_4697_5461# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X169 a_4701_3311# a_4535_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X170 VGND a_5843_4667# counter\[0\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X171 VPWR a_2971_8751# _026_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X172 a_6987_2197# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X173 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X174 VGND a_9586_6549# a_9515_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X175 VPWR a_8390_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X176 a_7323_4765# a_6541_4399# a_7239_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X177 VGND _004_ a_9933_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X179 VPWR _023_ a_1867_3561# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.265 ps=2.53 w=1 l=0.15
X180 a_7282_4221# counter\[0\] a_7193_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X181 VPWR counter\[5\] a_4771_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X182 VPWR _008_ a_7357_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X183 VGND _075_ a_2668_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X184 a_6719_10615# a_6887_10615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X185 VPWR a_2555_10704# a_2191_10615# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X186 VGND counter\[2\] a_7388_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X187 VGND net14 _028_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X189 a_1584_6351# _043_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X190 a_1827_6549# a_2111_6549# a_2046_6575# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X191 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X192 a_4227_2197# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X193 a_10287_6250# _082_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X194 a_5785_9813# counter\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X195 a_7745_7485# net10 a_7663_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X196 a_3601_2767# _014_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X197 a_3956_6391# _060_ a_3884_6391# VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X198 VGND _013_ a_4781_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X199 VGND net5 _024_ VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X200 VGND a_7171_10601# a_7178_10505# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X201 ones[8] a_9687_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X202 VPWR _084_ a_4627_5056# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X203 VPWR _061_ a_4627_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X204 VGND _073_ a_9503_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X205 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X206 _064_ a_3983_5056# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X207 VPWR a_4981_9991# _023_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X208 VGND a_7378_10660# a_7307_10761# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X209 a_5399_3677# a_4535_3311# a_5142_3423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X210 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X211 a_9629_9001# _087_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X212 ones[3] a_10239_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X213 a_7106_10749# a_6719_10615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X214 _058_ a_1867_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X215 VPWR net5 a_3123_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X216 VPWR counter\[8\] a_1683_10496# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X217 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X218 VGND a_2823_4943# a_2991_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X219 clknet_1_1__leaf_clk a_8390_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X220 a_6887_10615# a_7178_10505# a_7129_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X221 net14 a_7867_9019# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X222 VGND _090_ a_9624_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X223 VGND a_4215_4087# net13 VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X224 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X225 _010_ a_9435_9001# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X226 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X227 VPWR _060_ a_5363_2880# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X228 VGND a_6803_9813# a_6810_10113# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X229 net7 a_4279_2741# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X230 VPWR a_4123_9514# _009_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X231 a_6982_6005# a_6814_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X232 a_10287_6250# _082_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X233 a_4434_2197# a_4227_2197# a_4610_2589# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X234 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X236 clknet_1_0__leaf_clk a_4697_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X237 a_3295_10615# a_3391_10615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X238 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X239 VPWR _037_ a_4535_7232# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X240 VPWR clknet_1_0__leaf_clk a_6467_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X241 VGND _061_ a_4627_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X242 a_3701_5309# a_3431_4943# a_3611_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X243 VPWR a_5687_5175# _070_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X244 VGND _020_ a_5149_4233# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X245 VPWR _035_ a_4307_8439# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.074375 ps=0.815 w=0.42 l=0.15
X246 a_9899_4943# a_9117_4949# a_9815_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X247 VPWR net11 a_7847_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X248 a_4583_2223# a_4363_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X249 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X250 a_2129_7119# _017_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X251 VPWR a_5567_3579# a_5483_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X252 a_4610_2589# a_4363_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X253 VGND a_2191_10615# _056_ VGND sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X254 a_5250_4765# a_4977_4399# a_5165_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X255 a_9095_6549# a_9379_6549# a_9314_6575# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X256 a_5142_3423# a_4974_3677# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X257 _019_ a_6007_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X258 VPWR a_8447_8916# _006_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X259 VPWR a_9379_5461# a_9386_5761# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X260 VPWR a_7239_6031# a_7407_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X261 a_2111_6549# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X262 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X263 a_9687_4399# _049_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X264 a_4750_7913# _074_ a_4668_7913# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X265 VPWR a_8447_8439# _029_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X266 a_1460_9269# _059_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X267 a_5537_9839# counter\[9\] _090_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X268 VGND a_6169_6549# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X269 VPWR a_5675_4765# a_5843_4667# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X270 VGND a_4697_5461# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X271 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X272 VGND net14 a_10147_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X273 ones[1] a_9963_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X274 VGND _040_ a_5261_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X275 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X276 a_9739_6005# a_9915_6337# a_9867_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X277 VPWR a_4697_5461# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X278 a_4889_3311# _021_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X280 VPWR net7 a_7663_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X281 a_1581_5309# counter\[5\] a_1499_5056# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X282 VGND _054_ a_5087_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X283 VGND a_7791_9295# a_7959_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X284 a_2971_8751# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X285 VGND net8 a_2077_7691# VGND sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X287 a_7980_4649# _026_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X288 a_6607_2375# a_6703_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X289 a_3943_2197# a_4234_2497# a_4185_2589# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X290 _050_ _039_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X291 a_7123_2223# a_6987_2197# a_6703_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X292 VPWR clknet_1_0__leaf_clk a_4535_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X293 a_9091_8439# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X294 a_2313_4943# _018_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X295 VPWR _060_ a_3611_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X296 a_6003_10089# counter\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X297 VGND a_5675_4765# a_5843_4667# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X298 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X299 VPWR a_9213_3463# _063_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X300 clknet_0_clk a_6169_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X301 a_9841_4399# _049_ a_9769_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X302 clknet_1_0__leaf_clk a_4697_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X303 a_9091_8439# _060_ a_9325_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X304 VGND a_8447_8916# _006_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X305 VGND net1 a_4981_9991# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X306 a_6541_4399# a_6375_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X307 a_3295_10615# a_3391_10615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X308 VPWR a_3847_8903# _089_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X309 a_6173_3311# a_6007_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X310 VGND _080_ a_10045_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X311 a_4434_2197# a_4234_2497# a_4583_2223# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X312 a_7274_9117# a_6835_8751# a_7189_8751# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X314 a_9390_4943# a_8951_4949# a_9305_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X315 a_2111_6549# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X316 VPWR a_4279_2741# a_4195_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X317 VPWR a_8175_6549# _053_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X318 VGND _039_ a_8109_5639# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X319 a_4160_7479# a_3973_7119# a_4073_7235# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X320 a_1670_6351# net12 a_1584_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X321 a_8194_3561# _033_ a_7886_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X322 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X323 a_2191_10615# counter\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X325 VGND _009_ a_2665_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X326 _076_ a_2509_4663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X327 VPWR a_9091_10004# _002_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X328 a_9026_6031# a_8779_6409# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X329 a_6423_9991# a_6519_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X330 ones[8] a_9687_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X331 a_1941_7125# a_1775_7125# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X332 a_4771_2741# counter\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.31245 ps=1.68 w=0.42 l=0.15
X333 VPWR _036_ a_2879_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X334 a_4781_2223# a_4227_2197# a_4434_2197# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X335 VGND clknet_1_0__leaf_clk a_3247_2773# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X336 a_7400_8751# a_7001_8751# a_7274_9117# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X337 a_2509_4663# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X338 VPWR _072_ a_3799_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X339 a_9516_5321# a_9117_4949# a_9390_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X340 VPWR _090_ a_9896_9001# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X342 a_9205_4233# a_8215_3861# a_9079_3855# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X343 VGND a_8447_5175# _048_ VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X344 VPWR a_9815_4943# a_9983_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X345 VPWR a_8390_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X346 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X347 a_7171_10601# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X348 a_3029_6031# net6 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X349 VGND a_8631_2986# _014_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X350 _043_ a_7847_3133# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X351 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X352 VGND a_6719_10615# counter\[2\] VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X353 a_2214_7119# a_1775_7125# a_2129_7119# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X354 a_7357_9839# a_6810_10113# a_7010_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X355 VGND a_4595_4073# a_4602_3977# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X356 a_4311_4087# a_4602_3977# a_4553_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X357 VGND a_4697_5461# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X358 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X359 VGND counter\[2\] a_8209_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X360 ones[6] a_7939_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X361 a_2866_3087# net8 a_2697_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X362 a_9533_8751# counter\[10\] a_9624_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X363 VGND a_4123_9514# _009_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X364 VPWR a_7074_5599# a_7001_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X365 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X366 VGND a_9739_6005# _054_ VGND sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X367 _040_ a_4535_7232# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X368 VGND _063_ a_4137_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X369 a_9117_4949# a_8951_4949# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X370 a_2340_7497# a_1941_7125# a_2214_7119# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X371 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X372 a_2467_6575# a_2247_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X373 a_2723_7119# a_1941_7125# a_2639_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X375 a_2555_10704# counter\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X377 a_6887_10615# a_7171_10601# a_7106_10749# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X378 VPWR net7 a_9919_4087# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X379 VPWR _068_ a_5960_5175# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1087 ps=1.36 w=0.42 l=0.15
X380 a_6614_3423# a_6446_3677# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X381 a_9915_6337# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X382 a_6614_3423# a_6446_3677# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X383 VGND a_4802_4132# a_4731_4233# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X384 _041_ _028_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X385 a_10055_8527# counter\[0\] a_9961_8527# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X386 a_6982_4511# a_6814_4765# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X387 a_7274_9117# a_7001_8751# a_7189_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X389 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X390 a_8999_6727# a_9095_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X391 a_2542_3971# _086_ a_2460_3971# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X392 a_7917_9673# a_6927_9301# a_7791_9295# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X393 clknet_1_1__leaf_clk a_8390_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X394 net8 a_9247_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X395 VPWR clknet_1_0__leaf_clk a_1775_7125# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X396 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X397 VPWR a_10199_3285# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X398 _045_ a_4073_7235# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X399 ones[6] a_7939_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X400 a_4668_7913# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X401 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X402 clknet_0_clk a_6169_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X403 VPWR _060_ a_4627_5056# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X404 VPWR a_8263_6263# counter\[10\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X405 ones[1] a_9963_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X406 VGND a_7239_6031# a_7407_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X407 VGND _043_ a_8665_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X408 VGND a_7407_6005# a_7365_6409# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X409 VPWR a_8390_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X410 VGND a_10199_2197# net2 VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X411 a_9739_6005# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X412 a_7565_3311# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X413 clknet_1_0__leaf_clk a_4697_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X414 VPWR _039_ a_2409_9001# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X415 a_8850_6308# a_8650_6153# a_8999_6397# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X416 VPWR a_6423_9991# counter\[8\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X417 a_3983_5056# _062_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X418 VPWR a_6719_10615# counter\[2\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X419 VPWR _013_ a_4781_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X421 VPWR net1 a_2971_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X422 a_6761_10205# a_6423_9991# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X423 a_2398_4943# a_2125_4949# a_2313_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X424 _074_ a_1499_5056# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X425 clknet_0_clk a_6169_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X426 VPWR _074_ a_2513_3561# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X427 a_4457_8567# _028_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.122275 ps=1.08 w=0.42 l=0.15
X428 VGND a_8390_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X429 VPWR counter\[4\] a_5359_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X430 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X431 a_6423_9991# a_6519_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X432 ones[2] a_9871_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X433 VPWR clknet_1_1__leaf_clk a_8215_3861# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X434 VPWR a_7442_8863# a_7369_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X435 a_7281_9295# _012_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X436 a_4363_2223# a_4234_2497# a_3943_2197# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X437 VGND a_6169_6549# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X438 a_3675_10601# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X439 a_8076_3311# net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X440 a_9197_6409# a_8643_6249# a_8850_6308# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X441 a_9379_6549# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X442 a_2309_7119# a_1775_7125# a_2214_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X443 counter\[2\] a_6719_10615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X444 VGND a_4697_5461# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X445 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X446 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X447 a_7239_4765# a_6375_4399# a_6982_4511# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X448 clknet_1_1__leaf_clk a_8390_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X449 VPWR _023_ a_4535_7232# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X450 a_2318_6549# a_2118_6849# a_2467_6575# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X451 VPWR _048_ a_6007_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X452 VPWR _066_ a_5363_2880# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X453 VGND a_7111_4221# _068_ VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X454 a_7001_8751# a_6835_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X455 _092_ net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X456 a_9735_6575# a_9515_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X457 VPWR a_1731_6727# counter\[9\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X458 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X459 a_5418_4511# a_5250_4765# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X460 a_4617_7485# _023_ a_4535_7232# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X461 _035_ a_2866_3087# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X462 VGND net13 a_1670_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X463 VGND _043_ a_8657_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X464 a_10039_3087# net13 _050_ VGND sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X465 a_2021_4399# _056_ a_1949_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X466 a_2318_6549# a_2111_6549# a_2494_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X467 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X468 _060_ a_1460_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X469 a_8999_6727# a_9095_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X470 VGND net11 a_7847_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X471 a_2665_6575# a_2111_6549# a_2318_6549# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X472 _080_ a_3187_2251# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X473 VPWR _068_ a_3187_2251# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X474 a_9096_4373# net3 a_9319_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X475 VPWR a_2566_4917# a_2493_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X476 a_7111_4221# counter\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X477 a_6425_10602# _045_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X478 a_2494_6941# a_2247_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X479 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X480 a_8459_4551# net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X481 VPWR counter\[6\] _078_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X482 VPWR _050_ a_2787_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.265 ps=2.53 w=1 l=0.15
X483 a_8681_5309# _046_ a_8609_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X484 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X485 VPWR a_4521_8903# _025_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X486 a_8822_3829# a_8654_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X487 VGND _042_ a_8123_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X488 a_6391_2767# net2 _028_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X489 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X491 a_8459_4551# net11 a_8633_4427# VGND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X492 VPWR a_7407_4667# a_7323_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X494 a_2493_4943# a_1959_4949# a_2398_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X495 _073_ a_3799_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X496 _050_ net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X497 a_5149_4233# a_4602_3977# a_4802_4132# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X498 a_4521_8903# net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X499 a_8822_3829# a_8654_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X500 a_3882_10660# a_3682_10505# a_4031_10749# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X501 a_6922_2223# a_6607_2375# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X502 VPWR _004_ a_9933_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X503 _016_ a_7886_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X504 a_9379_6549# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X505 VPWR a_8459_4551# _042_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X506 a_9867_6397# _058_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X507 a_4889_3311# _021_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X508 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X509 a_5675_4765# a_4811_4399# a_5418_4511# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X510 VPWR _031_ a_8215_10496# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X511 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X512 VPWR a_5717_4087# _083_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X514 a_10199_3285# pulse VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X515 VPWR clknet_1_0__leaf_clk a_1959_4949# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X516 VGND a_5507_10357# _034_ VGND sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X517 a_3142_8751# net5 a_3053_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.06195 ps=0.715 w=0.42 l=0.15
X518 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X519 a_9586_6549# a_9386_6849# a_9735_6575# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X520 a_2665_6575# a_2118_6849# a_2318_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X521 VGND a_10195_7338# _020_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X522 VGND net1 a_3248_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.0693 ps=0.75 w=0.42 l=0.15
X523 VGND a_3882_10660# a_3811_10761# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X524 VPWR counter\[0\] _062_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X525 a_1653_5309# counter\[4\] a_1581_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X526 a_6906_5853# a_6467_5487# a_6821_5487# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X527 VGND a_6169_6549# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X528 VGND a_1731_6727# counter\[9\] VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X529 a_4345_6031# _091_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X530 _071_ counter\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X531 net4 a_5567_3579# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X532 _031_ _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X533 a_3610_10749# a_3295_10615# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X535 VPWR a_3675_10601# a_3682_10505# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X536 VGND a_6425_10602# _018_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X537 a_7554_10383# a_7307_10761# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X539 _051_ a_9687_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X540 VPWR clknet_1_0__leaf_clk a_6375_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X541 VPWR a_4697_5461# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X542 a_9586_6549# a_9379_6549# a_9762_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X543 a_4709_6825# _058_ _059_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X544 a_4731_4233# a_4602_3977# a_4311_4087# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X545 VPWR _037_ a_7663_7485# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X546 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X547 a_9933_6575# a_9379_6549# a_9586_6549# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X548 _026_ a_2971_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X549 VPWR net7 a_5507_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X551 a_7541_2223# a_6994_2497# a_7194_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X552 VPWR a_5843_4667# a_5759_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X553 _087_ a_7419_5281# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X555 _017_ _041_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X556 a_6738_9839# a_6423_9991# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X557 a_7378_10660# a_7171_10601# a_7554_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X558 a_1683_10496# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X559 a_9762_6941# a_9515_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X560 a_9095_5461# a_9386_5761# a_9337_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X561 a_9305_4943# _016_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X562 a_10045_10927# counter\[8\] _084_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X563 VPWR a_7407_6005# counter\[1\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X564 VPWR _068_ a_1683_10496# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X565 VGND a_7039_3579# a_6997_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X566 a_9595_3087# net11 a_9845_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X567 a_7388_4221# counter\[3\] a_7282_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X568 VGND _036_ a_2879_3855# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X569 a_8272_5737# net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X570 _065_ counter\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X571 _038_ a_6475_7913# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X572 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X573 VPWR a_6169_6549# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X574 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X575 a_7366_9295# a_7093_9301# a_7281_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X576 a_2513_3561# counter\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X577 ones[2] a_9871_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X578 a_1867_4399# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X579 VGND a_8109_5639# _044_ VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X580 a_2247_6575# a_2118_6849# a_1827_6549# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X581 clknet_1_1__leaf_clk a_8390_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X582 a_4232_7479# _028_ a_4160_7479# VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X583 a_1679_10089# _042_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X584 a_5359_4943# _068_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X585 clknet_0_clk a_6169_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X586 a_1679_10089# net12 a_1461_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X587 a_5149_4233# a_4595_4073# a_4802_4132# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X588 a_2787_8207# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1475 ps=1.295 w=1 l=0.15
X589 a_6729_6031# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X590 _067_ a_5363_2880# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X591 VPWR _027_ a_8447_8439# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.074375 ps=0.815 w=0.42 l=0.15
X592 a_7442_8863# a_7274_9117# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X593 a_7307_10761# a_7178_10505# a_6887_10615# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X594 VGND a_9815_4943# a_9983_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X595 VPWR a_8390_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X596 VPWR net10 a_5369_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X597 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X598 a_5717_4087# counter\[8\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X599 a_5517_3133# _065_ a_5445_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X600 VPWR net12 _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.135 ps=1.27 w=1 l=0.15
X601 a_9314_6575# a_8999_6727# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X602 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X603 clknet_1_0__leaf_clk a_4697_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X604 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X605 VPWR a_4434_2197# a_4363_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X606 _077_ a_4668_7913# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X607 a_9515_5487# a_9386_5761# a_9095_5461# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X608 a_5185_7913# _092_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X609 a_4431_6351# net3 _092_ VGND sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X610 a_5918_5303# _069_ a_5837_5303# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.05355 ps=0.675 w=0.42 l=0.15
X611 a_10039_3087# net12 a_9845_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X612 a_7331_5853# a_6467_5487# a_7074_5599# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X613 VPWR a_9919_4087# _033_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X614 VGND a_4279_2741# a_4237_3145# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X615 a_4771_2741# counter\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X616 VGND a_8263_6263# counter\[10\] VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X617 a_7825_8751# a_6835_8751# a_7699_9117# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X618 VPWR clknet_1_0__leaf_clk a_4811_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X619 VPWR _060_ a_9435_9001# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X620 _085_ a_4627_5056# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X621 a_9933_6575# a_9386_6849# a_9586_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X622 a_5507_10357# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.31245 ps=1.68 w=0.42 l=0.15
X623 a_4538_8567# _035_ a_4457_8567# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.05355 ps=0.675 w=0.42 l=0.15
X624 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X625 VGND a_8390_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X626 VGND _053_ _021_ VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X627 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X628 VPWR a_6515_4074# _013_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X629 VGND a_7867_9019# a_7825_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X630 VPWR a_7534_9269# a_7461_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X631 VPWR a_6871_3677# a_7039_3579# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X632 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X633 VPWR net4 _052_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X634 a_9941_5321# a_8951_4949# a_9815_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X635 net2 a_10199_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X636 a_6169_6549# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X637 a_7365_6409# a_6375_6037# a_7239_6031# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X638 _082_ a_3797_6147# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X639 VPWR a_8999_5639# counter\[4\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X640 VGND a_2566_4917# a_2524_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X641 VPWR a_7499_5755# a_7415_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X642 a_6283_7669# _037_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X643 _004_ a_9503_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X644 VPWR net13 a_10239_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X645 a_7461_9295# a_6927_9301# a_7366_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X646 ones[9] a_10239_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X647 VGND a_8643_6249# a_8650_6153# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X648 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X649 a_2765_7497# a_1775_7125# a_2639_7119# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X650 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X651 net8 a_9247_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X652 net3 a_7407_4667# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X653 clknet_1_0__leaf_clk a_4697_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X654 VPWR _069_ a_5687_5175# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.074375 ps=0.815 w=0.42 l=0.15
X655 a_8477_6575# net4 a_8175_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X656 a_7929_3133# net7 a_7847_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X657 a_2409_4445# _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X658 a_7505_5281# counter\[9\] a_7419_5281# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X659 ones[5] a_10239_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X660 VPWR net14 a_10147_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X663 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X664 a_2639_7119# a_1775_7125# a_2382_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X665 a_7699_9117# a_6835_8751# a_7442_8863# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X666 VPWR a_5785_9813# _066_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X667 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X668 VGND a_6607_2375# counter\[6\] VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X669 VPWR a_6169_6549# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X670 VPWR net3 a_10239_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X671 _091_ net14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X672 VPWR _009_ a_2665_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X673 ones[0] a_10239_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X674 VPWR _060_ a_3847_8903# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.074375 ps=0.815 w=0.42 l=0.15
X675 a_10081_4221# _026_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X676 a_4031_10749# a_3811_10761# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X677 VGND _007_ a_9933_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X678 clknet_0_clk a_6169_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X679 a_6519_9813# a_6803_9813# a_6738_9839# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X680 a_3675_10601# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X681 VGND a_7194_2197# a_7123_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X682 net3 a_7407_4667# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X683 a_5687_5175# _059_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.142225 ps=1.335 w=0.42 l=0.15
X684 VPWR a_7378_10660# a_7307_10761# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X685 a_7191_7119# _025_ _012_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.26 ps=2.52 w=1 l=0.15
X686 ones[0] a_10239_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X687 a_2313_4943# _018_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X689 a_1950_3311# _023_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.17225 ps=1.83 w=0.65 l=0.15
X690 a_9091_10004# _067_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X692 VGND a_6871_3677# a_7039_3579# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X693 VGND net13 a_10239_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X694 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X695 a_4974_3677# a_4535_3311# a_4889_3311# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X696 a_7093_9301# a_6927_9301# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X697 a_3882_10660# a_3675_10601# a_4058_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X698 ones[9] a_10239_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X699 VPWR counter\[5\] a_1499_5056# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X700 a_3854_2741# a_3686_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X701 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X702 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X703 a_9079_3855# a_8215_3861# a_8822_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X704 VPWR _055_ a_1867_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X705 VPWR a_4111_2767# a_4279_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X706 a_7290_7119# _024_ a_7191_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1725 ps=1.345 w=1 l=0.15
X707 a_4781_5309# _083_ a_4709_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X708 VPWR a_7867_9019# a_7783_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X709 VGND a_8999_5639# counter\[4\] VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X710 VPWR a_2807_7093# a_2723_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X711 ones[5] a_10239_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X712 a_7663_7485# net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X714 a_2682_3311# counter\[7\] a_2513_3561# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X716 a_4689_7485# _034_ a_4617_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X717 a_9961_8207# counter\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X718 clknet_0_clk a_6169_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X719 a_5507_10357# net6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X720 a_4229_10761# a_3675_10601# a_3882_10660# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X721 a_9595_3087# _039_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X722 VGND a_8390_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X723 VGND a_7407_6005# counter\[1\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X724 VGND a_9091_8439# _079_ VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X725 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X726 VGND clknet_1_0__leaf_clk a_6467_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X727 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X728 a_5399_3677# a_4701_3311# a_5142_3423# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X729 clknet_1_1__leaf_clk a_8390_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X730 _031_ net7 a_5541_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X731 a_4111_2767# a_3247_2773# a_3854_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X732 VGND counter\[9\] a_2460_3971# VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X736 VPWR _028_ a_7886_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X737 VPWR a_1461_9813# _047_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X738 VPWR a_9558_4917# a_9485_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X739 VPWR a_9247_3829# a_9163_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X740 a_8447_5175# _028_ a_8681_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X741 VGND a_9379_5461# a_9386_5761# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X743 VPWR a_3847_2375# net6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X744 VGND a_7867_9019# net14 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X745 _088_ a_2460_3971# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X746 a_6541_6037# a_6375_6037# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X747 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X748 clknet_1_1__leaf_clk a_8390_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X749 a_6987_2197# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X750 VPWR a_9832_8181# _069_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X751 VPWR net5 a_2971_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X752 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X753 VGND net2 _059_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X754 VGND clknet_1_1__leaf_clk a_8215_3861# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X755 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X756 a_9485_4943# a_8951_4949# a_9390_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X757 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X758 a_8393_6825# net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X759 VPWR a_9586_5461# a_9515_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X760 VPWR clk a_6169_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X761 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X762 VGND a_3675_10601# a_3682_10505# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X763 VPWR _050_ a_9687_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X764 VPWR a_4227_2197# a_4234_2497# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X765 VPWR counter\[2\] a_2191_10615# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X766 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X767 VGND a_8850_6308# a_8779_6409# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X768 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X769 a_9961_8207# counter\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X770 _061_ a_3611_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X771 VGND clknet_0_clk a_4697_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X772 clknet_1_0__leaf_clk a_4697_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X773 VPWR net8 a_1991_7691# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X774 a_8597_8567# _028_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.122275 ps=1.08 w=0.42 l=0.15
X775 VGND a_9096_4373# _093_ VGND sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X776 a_6909_6031# a_6375_6037# a_6814_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X778 net12 a_7499_5755# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X779 VGND a_4697_5461# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X780 VPWR clknet_1_1__leaf_clk a_8951_4949# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X781 a_4307_8439# _028_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.142225 ps=1.335 w=0.42 l=0.15
X782 VPWR counter\[4\] a_8338_11177# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X783 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X784 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X785 a_6871_3677# a_6007_3311# a_6614_3423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X786 a_8447_8916# _079_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X787 a_6391_2767# net14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X788 a_3686_2767# a_3247_2773# a_3601_2767# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X789 VPWR a_7867_9019# net14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X791 a_6169_6549# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X792 a_9225_4399# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X793 a_3847_8903# a_4120_8731# a_4078_8757# VGND sky130_fd_pr__nfet_01v8 ad=0.107825 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X794 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X795 VGND a_9213_3463# _063_ VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X796 VGND a_6169_6549# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X797 _086_ a_1683_10496# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X798 VPWR clknet_1_1__leaf_clk a_6375_6037# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X799 VGND clknet_1_1__leaf_clk a_6927_9301# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X801 net12 a_7499_5755# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X802 a_8109_5639# _039_ a_8272_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X803 a_7419_5281# counter\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X804 a_3812_3145# a_3413_2773# a_3686_2767# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X805 clknet_1_0__leaf_clk a_4697_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X806 VGND a_5142_3423# a_5100_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X807 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X808 a_8359_6263# a_8650_6153# a_8601_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X809 a_6814_4765# a_6375_4399# a_6729_4399# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X810 _037_ a_1991_7691# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X811 a_2214_7119# a_1941_7125# a_2129_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X812 VGND _033_ a_8076_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X813 VPWR a_2111_6549# a_2118_6849# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X814 VPWR a_6169_6549# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X815 _068_ a_7111_4221# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X816 VGND _066_ a_5517_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X817 VGND clknet_1_0__leaf_clk a_1959_4949# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X818 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X819 _011_ _093_ a_5185_7913# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X820 a_6803_9813# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X821 VGND a_6515_4074# _013_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X822 a_8447_8916# _079_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X823 a_8657_6575# net12 a_8561_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X824 counter\[0\] a_5843_4667# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X825 a_5507_10357# net7 a_5905_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X826 a_4111_2767# a_3413_2773# a_3854_2741# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X827 VGND _068_ a_6733_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X828 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X829 a_6940_4399# a_6541_4399# a_6814_4765# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X830 a_6423_11079# counter\[10\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X831 a_9319_4399# _091_ a_9225_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X832 a_1867_3561# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1475 ps=1.295 w=1 l=0.15
X833 _030_ a_7980_4649# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X834 a_6729_4399# _011_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X835 VGND clknet_0_clk a_8390_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X836 a_3973_7119# _043_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X837 a_7239_4765# a_6541_4399# a_6982_4511# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X838 VGND _026_ a_8720_8439# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10785 ps=1.36 w=0.42 l=0.15
X839 net5 a_7959_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X841 VGND net7 a_7980_4649# VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X842 VGND a_5141_4917# _075_ VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X843 VGND a_1461_9813# _047_ VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X845 a_3315_6351# net3 a_3219_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X846 VGND a_7699_9117# a_7867_9019# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X847 VPWR a_3973_7119# a_4073_7235# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X848 VPWR a_2382_7093# a_2309_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X849 VGND clknet_1_0__leaf_clk a_4535_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X850 counter\[0\] a_5843_4667# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X851 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X852 VPWR a_7959_9269# a_7875_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X853 VPWR _043_ a_1501_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X854 a_3811_10761# a_3675_10601# a_3391_10615# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X855 a_7111_4221# counter\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X856 _003_ a_2603_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X857 a_4802_4132# a_4595_4073# a_4978_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X858 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X859 a_8393_6825# _025_ a_8175_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X860 _072_ a_8256_11177# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X861 VGND a_9558_4917# a_9516_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X862 VPWR counter\[10\] _090_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X863 a_6173_3311# a_6007_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X864 VPWR a_6987_2197# a_6994_2497# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X865 VGND a_2111_6549# a_2118_6849# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X866 a_5703_10749# net3 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196275 ps=1.33 w=0.42 l=0.15
X867 a_7886_3311# _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X868 VGND _047_ sky130_fd_pr__diode_pw2nd_05v5 perim=2.64e+06 area=4.347e+11
X869 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X870 a_8850_6308# a_8643_6249# a_9026_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X871 VGND _072_ a_3953_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X872 a_9435_9001# counter\[10\] a_9629_9001# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X873 VGND a_10199_3285# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X874 a_2513_10749# counter\[3\] a_2413_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X875 a_7386_7439# net5 _012_ VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.115375 ps=1.005 w=0.65 l=0.15
X876 a_3811_10761# a_3682_10505# a_3391_10615# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X877 a_8907_2986# _085_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X878 VGND _006_ a_7541_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X879 a_9096_4373# net2 a_9225_4649# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X880 clknet_1_1__leaf_clk a_8390_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X881 a_3248_8751# net3 a_3142_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X882 a_2866_3087# _023_ a_2780_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X883 _028_ net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X884 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X885 VPWR a_6425_10602# _018_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X886 a_4697_5461# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X887 a_6088_9839# counter\[1\] a_5785_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X888 _073_ a_3799_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X889 VPWR a_4697_5461# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X890 a_10153_4221# net7 a_10081_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X891 VGND a_3295_10615# counter\[5\] VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X892 net4 a_5567_3579# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X893 VGND counter\[3\] a_9832_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X894 a_6423_11079# counter\[9\] a_6657_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X895 net9 a_9983_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X896 clknet_1_1__leaf_clk a_8390_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X897 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X898 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X899 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X901 VPWR net6 a_9871_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X902 a_5675_4765# a_4977_4399# a_5418_4511# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X903 VGND _023_ a_3315_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X904 a_9624_8751# _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X905 VPWR a_7699_9117# a_7867_9019# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X906 a_9921_3476# _076_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X907 VPWR a_6803_9813# a_6810_10113# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X908 VPWR clk a_6169_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X909 _003_ a_2603_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X910 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X911 clknet_0_clk a_6169_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X912 a_2596_3311# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X914 a_9305_4943# _016_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X915 a_5880_3971# counter\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X916 a_7194_2197# a_6987_2197# a_7370_2589# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X917 VPWR a_8390_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X918 VPWR counter\[6\] a_4750_7913# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X919 a_7001_8751# a_6835_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X920 VGND _084_ a_4781_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X921 clknet_1_0__leaf_clk a_4697_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X922 VPWR net12 a_9687_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X923 a_8678_8567# _027_ a_8597_8567# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.05355 ps=0.675 w=0.42 l=0.15
X924 _027_ a_3029_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X925 _032_ a_8215_10496# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X926 net10 a_2807_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X927 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X928 VPWR a_8447_5175# _048_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X929 a_9091_8439# _078_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X930 a_10195_7338# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X931 VGND a_4697_5461# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X932 VGND _081_ a_3956_6391# VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X934 ones[10] a_9687_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X935 a_7343_2223# a_7123_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X936 VGND _033_ a_4580_8439# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10785 ps=1.36 w=0.42 l=0.15
X937 a_7370_2589# a_7123_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X938 VGND a_6982_4511# a_6940_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X939 VGND _087_ a_4120_8731# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10785 ps=1.36 w=0.42 l=0.15
X940 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X941 VGND a_4307_8439# _036_ VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X942 a_9197_6409# a_8650_6153# a_8850_6308# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X943 a_8578_6397# a_8263_6263# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X944 a_4215_4087# a_4311_4087# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X945 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X946 clknet_0_clk a_6169_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X947 a_3847_2375# a_3943_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X948 VPWR _028_ a_9687_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X949 VGND a_8390_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X950 a_2191_10615# a_2555_10704# a_2513_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X951 a_3391_10615# a_3682_10505# a_3633_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X952 VPWR net10 a_7939_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X953 a_1827_6549# a_2118_6849# a_2069_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X954 VPWR a_7039_3579# a_6955_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X955 _080_ a_3187_2251# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X956 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X957 a_5141_4917# counter\[5\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X958 a_1461_9813# net12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X961 a_7129_10383# a_6719_10615# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X963 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X964 net11 a_2991_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X965 VGND _050_ a_9841_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X966 VGND net14 _091_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X967 VGND a_2382_7093# a_2340_7497# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X968 VPWR a_3295_10615# counter\[5\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X969 _078_ counter\[6\] a_7565_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X973 VPWR _007_ a_9933_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X974 a_8569_3855# _015_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X975 clknet_1_1__leaf_clk a_8390_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X976 VPWR a_4802_4132# a_4731_4233# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X977 a_2077_7691# net9 a_1991_7691# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X978 VGND a_2971_8751# _026_ VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X979 a_6703_2197# a_6994_2497# a_6945_2589# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X980 VGND counter\[0\] a_9213_3463# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X981 a_3797_6147# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X982 ones[10] a_9687_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X983 _016_ a_7886_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X984 VGND _048_ a_6007_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X985 a_4802_4132# a_4602_3977# a_4951_4221# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X986 a_8175_6549# _025_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X987 a_6821_5487# _019_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X988 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X989 a_7331_5853# a_6633_5487# a_7074_5599# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X990 VGND net10 a_7939_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X991 VGND a_9983_4917# a_9941_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X992 a_8643_6249# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X993 VGND clknet_1_0__leaf_clk a_6375_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X994 a_1501_6031# net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X995 VPWR counter\[2\] a_7111_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.0588 ps=0.7 w=0.42 l=0.15
X996 _049_ a_1670_6351# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X997 VPWR net5 a_9963_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X998 VPWR clknet_1_0__leaf_clk a_6007_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X999 _058_ a_1867_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1000 VGND a_5418_4511# a_5376_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1001 a_7194_2197# a_6994_2497# a_7343_2223# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1002 a_5250_4765# a_4811_4399# a_5165_4399# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1004 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1005 a_4981_9991# net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1006 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1007 VGND counter\[0\] a_9677_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1008 VPWR counter\[0\] a_3431_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1009 a_1731_6727# a_1827_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1010 a_3601_2767# _014_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1011 VGND clknet_0_clk a_8390_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1012 _039_ a_7663_7485# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X1013 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1014 _074_ a_1499_5056# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1015 _028_ net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1016 a_2382_7093# a_2214_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1017 a_3123_6031# net6 a_3029_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X1018 VPWR a_1460_9269# _060_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1019 a_7472_7439# net3 a_7386_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1020 VGND clknet_1_0__leaf_clk a_1775_7125# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1021 a_7541_2223# a_6987_2197# a_7194_2197# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1022 VGND clknet_0_clk a_4697_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1023 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1024 VGND counter\[0\] a_6088_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1025 a_3413_2773# a_3247_2773# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1026 a_5376_4399# a_4977_4399# a_5250_4765# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1027 clknet_1_0__leaf_clk a_4697_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1028 a_9095_6549# a_9386_6849# a_9337_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1029 a_6423_11079# counter\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1030 a_6939_9839# a_6810_10113# a_6519_9813# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1031 VPWR a_7331_5853# a_7499_5755# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1032 _010_ a_9435_9001# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1033 VPWR a_7111_4221# _068_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X1034 VGND net6 a_9871_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1035 VPWR counter\[7\] a_4771_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X1036 a_2413_10749# counter\[2\] a_2325_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X1037 a_9921_3476# _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1038 a_1949_4399# _055_ a_1867_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1039 VPWR _026_ a_7847_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1040 VPWR a_9739_6005# _054_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X1041 a_4595_4073# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1042 _035_ a_2866_3087# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1043 _046_ net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1044 a_8209_2223# counter\[0\] a_8113_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1045 a_3697_6031# _080_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1046 VPWR net13 _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0.135 ps=1.27 w=1 l=0.15
X1047 VGND net2 a_4521_8903# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1048 a_5165_4399# _000_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1049 a_3997_8757# _088_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.122275 ps=1.08 w=0.42 l=0.15
X1050 VGND a_6169_6549# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1051 a_2682_3311# counter\[6\] a_2596_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1052 a_4771_2741# counter\[5\] a_5169_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X1053 a_2566_4917# a_2398_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1054 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1055 VPWR _020_ a_5149_4233# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X1056 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1057 VPWR counter\[9\] a_2542_3971# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1058 VGND clknet_1_0__leaf_clk a_4811_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1059 VPWR a_6169_6549# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1060 clknet_1_1__leaf_clk a_8390_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1061 VGND a_2991_4917# a_2949_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1062 a_4981_9991# net1 a_5144_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1063 VGND net12 a_9687_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1064 VPWR _002_ a_7725_10761# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X1065 a_9515_6575# a_9386_6849# a_9095_6549# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1066 a_4697_5461# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1067 VGND _031_ a_6475_7913# VGND sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1068 VPWR a_4697_5461# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1069 a_5759_4765# a_4977_4399# a_5675_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1070 VPWR counter\[0\] a_9961_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1071 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1072 VGND _068_ a_1837_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1073 a_4974_3677# a_4701_3311# a_4889_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1074 a_9337_5853# a_8999_5639# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X1075 _060_ a_1460_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1076 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1077 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1078 VPWR _010_ a_9197_6409# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X1079 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1080 VGND clknet_1_1__leaf_clk a_8951_4949# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1081 VGND net2 a_9915_6337# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1082 a_4058_10383# a_3811_10761# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X1083 a_2566_4917# a_2398_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1084 net10 a_2807_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1085 a_1731_6727# a_1827_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1086 a_8631_2986# _032_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1087 VPWR a_9079_3855# a_9247_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1088 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1089 a_9253_8573# _078_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X1090 net1 a_10199_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1091 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1092 VGND a_7074_5599# a_7032_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1093 clknet_0_clk a_6169_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1094 VPWR a_8390_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1095 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1096 a_7442_8863# a_7274_9117# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1098 VPWR a_8999_6727# counter\[7\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1099 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1100 clknet_1_0__leaf_clk a_4697_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1101 net2 a_10199_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1102 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1103 a_8447_8439# _028_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.142225 ps=1.335 w=0.42 l=0.15
X1104 net5 a_7959_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1105 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1106 _022_ a_5087_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1107 a_8907_2986# _085_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1108 a_9515_5487# a_9379_5461# a_9095_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X1109 a_4530_4221# a_4215_4087# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X1110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1111 VPWR _006_ a_7541_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X1112 a_7032_5487# a_6633_5487# a_6906_5853# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1113 a_2823_4943# a_1959_4949# a_2566_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1114 a_9390_4943# a_9117_4949# a_9305_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1115 a_8447_5175# _028_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1116 VGND a_3847_8903# _089_ VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X1117 a_3391_10615# a_3675_10601# a_3610_10749# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1118 _076_ a_2509_4663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1119 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1120 a_3273_2251# _055_ a_3187_2251# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1121 a_4345_6031# net1 _092_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1122 a_1670_6351# net13 a_1501_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X1123 a_6557_7913# a_6283_7669# a_6475_7913# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1124 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1125 VGND a_4771_2741# _055_ VGND sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X1126 VGND net5 a_9963_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1127 a_8447_8439# a_8720_8439# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1085 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1128 net9 a_9983_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1129 VPWR clknet_1_1__leaf_clk a_6835_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1130 a_6814_6031# a_6541_6037# a_6729_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1132 VGND _080_ a_5717_4087# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1133 a_3686_2767# a_3413_2773# a_3601_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1134 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1135 VPWR a_9379_6549# a_9386_6849# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1136 _052_ net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1137 a_8390_7119# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1138 VPWR net11 _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X1139 a_9919_4087# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X1140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1141 VPWR a_2318_6549# a_2247_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X1142 VPWR a_4697_5461# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1143 a_7534_9269# a_7366_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1144 a_8263_6263# a_8359_6263# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1145 VGND net1 a_7472_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.089375 ps=0.925 w=0.65 l=0.15
X1146 VGND a_7010_9813# a_6939_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X1147 a_4977_4399# a_4811_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1148 a_4065_5309# _060_ a_3983_5056# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1149 a_7833_7485# net7 a_7745_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1150 VGND _044_ a_4232_7479# VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X1151 _011_ _092_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1152 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1153 VPWR a_2991_4917# a_2907_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1154 _000_ a_4627_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1155 _004_ a_9503_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1156 a_6729_4399# _011_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1157 a_5717_4087# _080_ a_5880_3971# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1158 VPWR _087_ a_4120_8731# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1087 ps=1.36 w=0.42 l=0.15
X1159 a_8749_3855# a_8215_3861# a_8654_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1160 VGND a_8999_6727# counter\[7\] VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1161 VGND _031_ a_8369_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1162 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1163 VGND a_4697_5461# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1164 VGND net8 a_10239_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1165 VGND a_7534_9269# a_7492_9673# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1166 ones[4] a_10239_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1167 VGND counter\[4\] a_8256_11177# VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1168 a_7847_3133# _037_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1169 a_8654_3855# a_8215_3861# a_8569_3855# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1170 VGND counter\[7\] a_2682_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X1171 VPWR a_6982_6005# a_6909_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1173 VPWR a_3854_2741# a_3781_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1174 a_9376_3561# counter\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X1175 _085_ a_4627_5056# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1176 VGND _068_ a_1653_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1177 VPWR _005_ a_4229_10761# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X1178 a_4123_9514# _089_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1179 a_8633_4427# net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X1180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1181 a_7534_9269# a_7366_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1182 clknet_0_clk a_6169_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1183 VPWR a_8390_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1185 a_2780_3087# _034_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1187 a_5687_5175# a_5960_5175# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1085 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1188 _000_ a_4627_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1189 VGND _086_ a_7505_5281# VGND sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1190 net11 a_2991_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1191 a_3781_2767# a_3247_2773# a_3686_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1192 VGND a_9379_6549# a_9386_6849# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1193 _001_ a_4903_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1194 a_8780_4233# a_8381_3861# a_8654_3855# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1195 ones[7] a_7847_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1196 a_5483_3677# a_4701_3311# a_5399_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1197 a_4237_3145# a_3247_2773# a_4111_2767# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1199 a_4967_3133# counter\[6\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196275 ps=1.33 w=0.42 l=0.15
X1200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1201 a_7976_3311# _028_ a_7886_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X1202 a_5363_2880# _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1203 _062_ counter\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1204 VPWR net2 a_4709_6825# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1206 VGND a_5399_3677# a_5567_3579# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1207 a_3847_8903# a_4120_8731# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1085 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1208 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1209 a_6519_9813# a_6810_10113# a_6761_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1211 VGND a_8175_6549# _053_ VGND sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X1212 a_9079_3855# a_8381_3861# a_8822_3829# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1213 a_4215_4087# a_4311_4087# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1214 VPWR a_9586_6549# a_9515_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X1215 a_7281_9295# _012_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1216 a_3219_6351# net5 a_3029_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1217 a_6803_9813# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1218 a_4307_8439# a_4580_8439# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1085 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1219 VPWR a_6169_6549# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1220 clknet_1_1__leaf_clk a_8390_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1221 ready a_10147_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1222 a_2823_4943# a_2125_4949# a_2566_4917# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1223 counter\[3\] a_7039_3579# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1224 a_10199_2197# rst VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1225 a_7725_10761# a_7178_10505# a_7378_10660# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X1226 VPWR a_4697_5461# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1227 clknet_1_1__leaf_clk a_8390_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1228 VGND a_4434_2197# a_4363_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X1229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1230 a_1499_5056# counter\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1232 a_6633_5487# a_6467_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1234 _081_ a_2682_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1235 a_8999_6397# a_8779_6409# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X1236 _022_ a_5087_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1237 a_9379_5461# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1238 VPWR net7 a_10239_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1240 a_4185_2589# a_3847_2375# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X1241 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1242 a_5905_10749# net6 a_5799_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X1243 a_8393_6825# _043_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1244 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1245 a_7791_9295# a_6927_9301# a_7534_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1246 counter\[1\] a_7407_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1247 a_9845_3087# net11 a_9595_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1249 VPWR net3 a_4345_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X1250 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1251 a_9225_4649# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1252 a_6729_6031# _001_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1254 a_5069_3677# a_4535_3311# a_4974_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1255 a_5687_5175# a_5960_5175# a_5918_5303# VGND sky130_fd_pr__nfet_01v8 ad=0.107825 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1256 a_5100_3311# a_4701_3311# a_4974_3677# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1257 a_8256_11177# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1258 VGND _060_ a_3701_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1259 VPWR counter\[8\] a_6423_11079# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X1260 VPWR _081_ a_3797_6147# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1261 VGND _057_ a_2021_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1262 VPWR a_7194_2197# a_7123_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X1263 a_7323_6031# a_6541_6037# a_7239_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1264 _072_ a_8256_11177# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1265 VGND a_8447_8439# _029_ VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X1266 a_4195_2767# a_3413_2773# a_4111_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1267 _021_ _053_ a_2787_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1268 a_8359_6263# a_8643_6249# a_8578_6397# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1269 a_6871_3677# a_6173_3311# a_6614_3423# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1270 _050_ net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X1271 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1272 a_3847_2375# a_3943_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1275 a_4363_2223# a_4227_2197# a_3943_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X1276 VPWR _070_ a_2603_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1277 VPWR _039_ _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1278 a_4701_3311# a_4535_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1279 a_8123_3133# _037_ a_8017_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1280 VGND a_4521_8903# _025_ VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1281 VGND a_5843_4667# a_5801_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1282 _064_ a_3983_5056# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1283 VPWR _042_ a_7847_3133# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1284 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1286 a_8631_2986# _032_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1287 clknet_1_0__leaf_clk a_4697_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1288 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1290 VPWR a_6423_11079# _057_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X1291 a_6821_5487# _019_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1292 a_4553_3855# a_4215_4087# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X1293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1294 a_3943_2197# a_4227_2197# a_4162_2223# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1295 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1296 a_9769_4399# _028_ a_9687_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1297 VPWR a_6169_6549# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1298 a_8390_7119# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1299 a_4227_2197# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1300 VPWR counter\[0\] a_7111_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.07455 ps=0.775 w=0.42 l=0.15
X1301 VGND a_9079_3855# a_9247_3829# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1302 VGND a_4227_2197# a_4234_2497# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1303 VPWR a_7239_4765# a_7407_4667# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1304 clknet_0_clk a_6169_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1306 a_8447_5175# _047_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X1307 a_4123_9514# _089_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1308 a_3881_10927# _060_ a_3799_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1309 VPWR a_7499_5755# net12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1310 _024_ net3 a_1950_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
X1311 VPWR a_2191_10615# _056_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1313 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1314 VGND a_5785_9813# _066_ VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1315 a_9558_4917# a_9390_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1316 a_3413_2773# a_3247_2773# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1317 a_7186_10205# a_6939_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X1318 VGND _070_ a_2603_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1319 VGND a_5687_5175# _070_ VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X1320 VPWR clknet_0_clk a_8390_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1321 _001_ a_4903_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1322 a_6955_3677# a_6173_3311# a_6871_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1323 a_6585_10927# counter\[10\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X1324 a_7193_4221# counter\[1\] a_7111_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.1092 ps=1.36 w=0.42 l=0.15
X1325 VPWR _063_ a_3983_5056# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1326 VGND _002_ a_7725_10761# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1327 VPWR _073_ a_9503_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1328 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1329 _061_ a_3611_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X1330 a_4595_4073# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1331 a_6909_4765# a_6375_4399# a_6814_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1332 _026_ a_2971_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.17515 ps=1.265 w=0.65 l=0.15
X1333 VGND a_7239_4765# a_7407_4667# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1334 a_4731_4233# a_4595_4073# a_4311_4087# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X1335 VGND a_4111_2767# a_4279_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1336 VGND a_7499_5755# net12 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1337 a_7010_9813# a_6803_9813# a_7186_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X1338 VPWR a_8109_5639# _044_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X1339 VPWR a_10287_6250# _007_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1340 VPWR net4 a_9687_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1341 VPWR _064_ a_4903_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1342 VPWR _086_ a_7419_5281# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1343 clknet_0_clk a_6169_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1344 VGND a_6982_6005# a_6940_6409# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1345 VGND a_2318_6549# a_2247_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X1346 a_6945_2589# a_6607_2375# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X1347 VPWR counter\[1\] _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1348 VGND _008_ a_7357_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1349 VGND a_8390_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1350 a_9919_4087# net8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1351 a_4684_9001# net14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X1352 a_7457_5487# a_6467_5487# a_7331_5853# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1353 a_8779_6409# a_8643_6249# a_8359_6263# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X1354 a_8076_3311# _038_ a_7976_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X1355 a_9815_4943# a_8951_4949# a_9558_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1356 a_5165_4399# _000_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1357 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1358 VGND _037_ a_4689_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1359 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1360 _077_ a_4668_7913# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X1361 VGND a_6614_3423# a_6572_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1362 VGND net7 a_10239_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1363 _040_ a_4535_7232# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1364 VPWR a_9091_8439# _079_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X1365 a_6446_3677# a_6007_3311# a_6361_3311# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1366 a_3431_4943# counter\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1367 VGND a_9586_5461# a_9515_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X1368 VGND a_7499_5755# a_7457_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1369 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1370 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1371 VPWR a_9921_3476# _005_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1372 VGND _039_ a_9595_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1373 a_3953_10927# _071_ a_3881_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1374 VGND a_8459_4551# _042_ VGND sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1375 a_4137_5309# _062_ a_4065_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1376 a_1941_7125# a_1775_7125# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1377 _086_ a_1683_10496# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1378 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1379 VGND a_9091_10004# _002_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1380 VPWR counter\[1\] a_6003_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1381 _024_ net5 a_1867_3561# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1382 VGND a_10287_6250# _007_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1383 clknet_1_1__leaf_clk a_8390_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1384 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1385 a_5261_7439# _028_ _041_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1387 a_6572_3311# a_6173_3311# a_6446_3677# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1388 a_4627_5056# _083_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1389 VPWR a_3882_10660# a_3811_10761# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X1390 a_8062_4649# _026_ a_7980_4649# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1391 a_8263_6263# a_8359_6263# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1392 a_9533_8751# _060_ a_9435_9001# VGND sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X1393 _019_ a_6007_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1394 counter\[1\] a_7407_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1395 a_4951_4221# a_4731_4233# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X1396 a_6657_10927# counter\[8\] a_6585_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1397 VGND net4 a_9687_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1398 a_5063_3133# counter\[7\] a_4967_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X1399 _045_ a_4073_7235# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X1400 _068_ a_7111_4221# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.27995 ps=1.615 w=1 l=0.15
X1401 a_7159_9839# a_6939_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X1402 VPWR a_9983_4917# a_9899_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1403 VGND a_9247_3829# a_9205_4233# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1404 VPWR a_6607_2375# counter\[6\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1405 a_5541_6575# _026_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1406 a_4073_7235# _028_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X1407 VGND clknet_1_1__leaf_clk a_6375_6037# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1408 a_2460_3971# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1409 VPWR _077_ a_9091_8439# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X1410 ones[7] a_7847_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1411 a_6361_3311# _003_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1413 _051_ a_9687_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1414 a_2409_9001# _041_ _017_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1416 VGND a_4697_5461# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1417 a_9213_3463# counter\[0\] a_9376_3561# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1418 clknet_1_0__leaf_clk a_4697_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1419 _059_ _058_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1420 _015_ a_2879_3855# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1421 a_8381_3861# a_8215_3861# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1422 VPWR net4 a_8393_6825# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1423 VPWR a_8850_6308# a_8779_6409# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X1424 a_1460_9269# _059_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1425 a_6906_5853# a_6633_5487# a_6821_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1426 VGND a_6987_2197# a_6994_2497# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1427 a_4535_7232# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1428 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1429 a_2129_7119# _017_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1430 VPWR a_5141_4917# _075_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1431 _043_ a_7847_3133# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X1432 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1433 clknet_0_clk a_6169_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1434 VPWR a_8390_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1435 a_2382_7093# a_2214_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1436 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1437 a_8109_5639# net11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1438 a_1991_7691# net9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1439 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1440 _038_ a_6475_7913# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X1441 VPWR _060_ a_3799_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1442 a_7847_3133# net7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X1443 a_6814_6031# a_6375_6037# a_6729_6031# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1444 VGND a_6169_6549# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1445 a_8297_10749# _028_ a_8215_10496# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1446 VGND net8 a_2866_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X1447 a_9095_5461# a_9379_5461# a_9314_5487# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1448 VPWR net11 a_8459_4551# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1449 a_2596_4405# a_2409_4445# a_2509_4663# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X1450 a_2325_10749# counter\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X1451 a_3611_4943# a_3431_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1452 VPWR a_2409_4445# a_2509_4663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X1453 a_7699_9117# a_7001_8751# a_7442_8863# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1454 VGND a_7959_9269# a_7917_9673# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1455 VGND _005_ a_4229_10761# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1456 a_2069_6941# a_1731_6727# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X1457 clknet_1_1__leaf_clk a_8390_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1459 clknet_1_0__leaf_clk a_4697_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1460 VPWR _057_ a_1867_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1461 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1462 a_6940_6409# a_6541_6037# a_6814_6031# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1463 a_10195_7338# _051_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1464 a_5799_10749# net5 a_5703_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X1465 VGND _068_ a_5960_5175# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10785 ps=1.36 w=0.42 l=0.15
X1466 a_7010_9813# a_6810_10113# a_7159_9839# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1467 VPWR net14 a_6391_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1468 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1469 a_2697_2767# _023_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1470 a_9815_4943# a_9117_4949# a_9558_4917# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1471 a_7378_10660# a_7178_10505# a_7527_10749# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1472 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1473 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1474 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1475 a_9624_8751# _087_ a_9533_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X1476 a_2191_10615# counter\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X1477 a_7239_6031# a_6541_6037# a_6982_6005# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1478 a_8609_5309# _047_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X1479 a_2870_8527# _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.17225 ps=1.83 w=0.65 l=0.15
X1480 VGND _064_ a_4903_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1481 VPWR _075_ a_2509_4663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1482 a_2125_4949# a_1959_4949# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1483 a_7001_5853# a_6467_5487# a_6906_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1484 VGND a_7331_5853# a_7499_5755# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1485 a_5142_3423# a_4974_3677# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1486 a_2639_7119# a_1941_7125# a_2382_7093# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1487 a_7357_9839# a_6803_9813# a_7010_9813# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1488 a_1765_10749# counter\[8\] a_1683_10496# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1489 a_6169_6549# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1490 VPWR clknet_0_clk a_8390_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1491 VPWR _068_ _071_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1492 VPWR net7 _031_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1494 a_7189_8751# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1495 a_2247_6575# a_2111_6549# a_1827_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X1496 a_7663_7485# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1497 VGND a_9921_3476# _005_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1498 a_3973_7119# _043_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1499 a_5525_3311# a_4535_3311# a_5399_3677# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1500 VPWR _026_ a_8720_8439# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1087 ps=1.36 w=0.42 l=0.15
X1501 a_8369_10749# _030_ a_8297_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1502 a_5444_5263# counter\[4\] a_5141_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1503 a_7939_7485# _026_ a_7833_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1504 a_1764_9839# _040_ a_1461_9813# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1505 a_6541_4399# a_6375_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1506 a_3123_6031# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X1507 VGND a_5567_3579# a_5525_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1508 VGND _091_ a_4431_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
X1509 a_8665_3311# net12 _046_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1510 a_6733_7439# counter\[4\] _071_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1511 _090_ counter\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1512 VGND a_8390_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1513 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1514 _032_ a_8215_10496# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1515 VPWR net8 a_10239_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1516 a_7239_6031# a_6375_6037# a_6982_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1517 ones[4] a_10239_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1518 VGND a_6169_6549# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1519 a_8654_3855# a_8381_3861# a_8569_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1520 a_4781_2223# a_4234_2497# a_4434_2197# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X1521 VPWR a_5418_4511# a_5345_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1522 a_9337_6941# a_8999_6727# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X1523 VGND _039_ _017_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1524 VPWR _060_ a_3983_5056# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1525 a_6939_9839# a_6803_9813# a_6519_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X1526 a_7123_2223# a_6994_2497# a_6703_2197# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1527 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1528 VPWR clknet_0_clk a_4697_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1529 a_5359_4943# counter\[5\] a_5141_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1530 VPWR a_9096_4373# _093_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1531 VPWR counter\[2\] _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1532 VGND a_6423_9991# counter\[8\] VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1533 a_9919_4087# net8 a_10153_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1534 a_5345_4765# a_4811_4399# a_5250_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1535 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1536 VPWR a_4697_5461# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1537 VGND a_7442_8863# a_7400_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1538 a_6515_4074# _029_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1539 a_4978_3855# a_4731_4233# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X1540 VGND clknet_1_0__leaf_clk a_6007_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1541 VPWR net5 a_7290_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1542 VPWR _044_ a_4073_7235# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1543 a_5144_10089# net14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X1544 a_1837_10749# _055_ a_1765_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1545 a_7415_5853# a_6633_5487# a_7331_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1546 a_9832_8181# counter\[3\] a_9961_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1547 a_9225_4649# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1548 VGND _037_ a_6283_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X1549 net1 a_10199_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1550 a_2971_8751# net6 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.1092 ps=1.36 w=0.42 l=0.15
X1551 VGND net2 _028_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1552 _021_ _052_ a_2870_8527# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
X1553 VPWR a_6169_6549# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1554 VPWR a_7407_6005# a_7323_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1555 VPWR a_8822_3829# a_8749_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1557 _050_ net13 a_10039_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1558 VPWR _023_ a_3123_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X1559 a_5369_7119# _040_ _041_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X1560 VPWR a_5399_3677# a_5567_3579# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1561 a_9515_6575# a_9379_6549# a_9095_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X1562 a_5261_7439# net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1563 clknet_0_clk a_6169_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1565 a_3187_2251# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1566 clknet_1_0__leaf_clk a_4697_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1567 a_9091_10004# _067_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1568 VPWR _080_ _084_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1569 a_8017_3133# _026_ a_7929_3133# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1570 VPWR a_5507_10357# _034_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X1571 ready a_10147_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1572 VGND a_8390_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1573 a_5445_3133# _060_ a_5363_2880# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1574 a_8999_5639# a_9095_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1575 _037_ a_1991_7691# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1576 VGND a_5717_4087# _083_ VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1577 counter\[3\] a_7039_3579# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1578 a_2949_5321# a_1959_4949# a_2823_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1579 VPWR net5 a_5507_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X1580 VPWR _043_ _046_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1581 VPWR a_10199_2197# net2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1582 _027_ a_3029_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X1583 a_8447_8439# a_8720_8439# a_8678_8567# VGND sky130_fd_pr__nfet_01v8 ad=0.107825 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1584 _078_ _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1585 a_7189_8751# _022_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1586 a_4521_8903# net2 a_4684_9001# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1587 _028_ net2 a_6391_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1588 VPWR a_7010_9813# a_6939_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X1589 VPWR _033_ a_4580_8439# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1087 ps=1.36 w=0.42 l=0.15
X1590 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1591 VPWR a_7407_4667# net3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1592 VGND clknet_1_1__leaf_clk a_6835_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1593 a_4977_4399# a_4811_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1594 VPWR net12 a_8393_6825# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1595 VPWR a_4307_8439# _036_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X1596 a_3847_8903# _088_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.142225 ps=1.335 w=0.42 l=0.15
X1597 VPWR a_9915_6337# a_9739_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1598 VPWR a_2639_7119# a_2807_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1599 a_8643_6249# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1600 _082_ a_3797_6147# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X1601 VGND a_1460_9269# _060_ VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1602 VPWR _091_ a_9225_4649# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1603 VPWR a_8907_2986# _008_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1604 a_8561_6575# net13 a_8477_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1605 clknet_1_1__leaf_clk a_8390_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1606 VPWR net9 a_8194_3561# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X1607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1608 VPWR a_4215_4087# net13 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1609 a_4162_2223# a_3847_2375# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X1610 VGND clk a_6169_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1611 a_8390_7119# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1612 VGND a_3847_2375# net6 VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1613 a_6982_4511# a_6814_4765# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1614 a_7783_9117# a_7001_8751# a_7699_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1615 _087_ a_7419_5281# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1616 a_6607_2375# a_6703_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1617 VPWR net7 a_8062_4649# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1618 a_3884_6391# a_3697_6031# a_3797_6147# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X1619 a_7527_10749# a_7307_10761# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X1620 a_6361_3311# _003_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1621 VGND a_7407_4667# net3 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1622 VPWR net14 _091_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1623 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1624 _015_ a_2879_3855# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1626 a_8779_6409# a_8650_6153# a_8359_6263# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1627 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1628 clknet_1_0__leaf_clk a_4697_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1629 a_6997_3311# a_6007_3311# a_6871_3677# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1630 a_9735_5487# a_9515_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X1631 a_7365_4399# a_6375_4399# a_7239_4765# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1632 _091_ net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1633 VGND _068_ a_5444_5263# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1634 VGND _042_ a_1764_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1635 VPWR _040_ a_1679_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1636 VPWR a_7171_10601# a_7178_10505# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1637 VPWR a_10195_7338# _020_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1638 a_7307_10761# a_7171_10601# a_6887_10615# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 ones[6] ones[2] 0.137271f
C1 _007_ net13 0.412636f
C2 _023_ _035_ 0.21814f
C3 net14 counter\[9\] 0.464051f
C4 _088_ _027_ 0.133536f
C5 _038_ _093_ 0.125836f
C6 _043_ _022_ 0.138557f
C7 a_4627_5056# _084_ 0.215652f
C8 ones[7] _084_ 1.31569f
C9 a_7847_3855# VPWR 0.233915f
C10 _088_ VPWR 0.650891f
C11 _058_ _004_ 0.112457f
C12 _086_ counter\[9\] 0.8346f
C13 ones[6] _010_ 0.296857f
C14 a_9247_3829# VPWR 0.380984f
C15 a_2191_10615# VPWR 0.357234f
C16 a_1941_7125# a_2382_7093# 0.110715f
C17 a_1775_7125# a_2214_7119# 0.273138f
C18 net7 net11 0.323319f
C19 _071_ counter\[1\] 0.132501f
C20 a_5960_5175# VPWR 0.16387f
C21 net7 _045_ 0.104779f
C22 net14 _067_ 0.13435f
C23 net5 counter\[9\] 0.110698f
C24 a_7331_5853# VPWR 0.176013f
C25 _033_ counter\[3\] 0.103536f
C26 counter\[0\] _068_ 0.283115f
C27 _074_ net9 0.541951f
C28 _000_ _060_ 0.16076f
C29 _058_ _074_ 0.291928f
C30 _016_ clknet_1_1__leaf_clk 0.144913f
C31 _069_ _004_ 0.219948f
C32 _025_ _039_ 0.217483f
C33 _048_ _026_ 0.152583f
C34 net5 _067_ 0.465529f
C35 a_7039_3579# VPWR 0.443585f
C36 a_4111_2767# VPWR 0.193801f
C37 clknet_1_0__leaf_clk _003_ 0.398317f
C38 counter\[4\] a_8256_11177# 0.172112f
C39 _061_ _060_ 0.224222f
C40 net5 a_2971_8751# 0.16256f
C41 _045_ net9 0.359744f
C42 _034_ _015_ 0.14161f
C43 _060_ _073_ 0.134817f
C44 _045_ _041_ 0.307914f
C45 net14 net3 0.401915f
C46 _030_ VPWR 0.968279f
C47 _022_ _026_ 0.241659f
C48 _028_ _027_ 1.37624f
C49 _086_ net3 0.439198f
C50 _005_ net6 0.112687f
C51 _028_ net4 1.3266f
C52 _037_ _026_ 0.646919f
C53 counter\[5\] _085_ 0.127431f
C54 _088_ _015_ 0.316114f
C55 net1 _001_ 0.479487f
C56 _014_ VPWR 0.761426f
C57 _028_ VPWR 3.36887f
C58 counter\[2\] _026_ 1.14042f
C59 _091_ VPWR 0.740566f
C60 _054_ net12 0.275485f
C61 a_5418_4511# a_5250_4765# 0.239923f
C62 net5 net3 1.87336f
C63 _068_ net10 0.36536f
C64 counter\[6\] _028_ 0.38099f
C65 a_6987_2197# counter\[0\] 0.114096f
C66 _074_ _056_ 0.233578f
C67 a_3943_2197# VPWR 0.191909f
C68 a_2409_4445# _074_ 0.140004f
C69 a_1461_9813# _047_ 0.161092f
C70 _048_ counter\[3\] 0.103343f
C71 _037_ a_1991_7691# 0.11001f
C72 a_6446_3677# a_6007_3311# 0.260055f
C73 _018_ VPWR 1.88156f
C74 a_5087_6575# _022_ 0.108099f
C75 a_7123_2223# VPWR 0.190502f
C76 a_8447_8439# VPWR 0.203289f
C77 counter\[0\] _087_ 0.18018f
C78 _020_ _011_ 0.103059f
C79 _003_ a_2603_10927# 0.12546f
C80 a_9558_4917# a_9390_4943# 0.239923f
C81 counter\[5\] a_2125_4949# 0.236442f
C82 a_8951_4949# _028_ 0.182801f
C83 _010_ counter\[1\] 0.163107f
C84 _037_ counter\[3\] 0.214427f
C85 clknet_1_0__leaf_clk _060_ 0.561115f
C86 counter\[2\] counter\[3\] 0.688098f
C87 _086_ _080_ 0.860401f
C88 net7 net2 0.156992f
C89 counter\[4\] _037_ 1.01326f
C90 _016_ _063_ 0.194469f
C91 net1 net12 0.132567f
C92 _028_ a_4307_8439# 0.223501f
C93 net1 _077_ 0.2617f
C94 net3 clknet_1_1__leaf_clk 0.335595f
C95 counter\[7\] _084_ 0.388511f
C96 net12 net13 0.450591f
C97 net3 _059_ 0.16077f
C98 _053_ _042_ 0.160188f
C99 _082_ VPWR 0.496235f
C100 a_1959_4949# a_2566_4917# 0.136009f
C101 clknet_1_0__leaf_clk _042_ 0.137014f
C102 _058_ net2 0.107712f
C103 a_1959_4949# counter\[4\] 0.453131f
C104 a_3675_10601# a_3682_10505# 0.973502f
C105 _032_ counter\[7\] 0.263532f
C106 _042_ a_8459_4551# 0.110214f
C107 ones[8] VPWR 0.262905f
C108 a_4697_5461# net11 0.136252f
C109 a_9117_4949# counter\[2\] 0.27408f
C110 _034_ _036_ 0.381512f
C111 a_8359_6263# a_8650_6153# 0.192261f
C112 _027_ VPWR 1.96606f
C113 _026_ _024_ 0.913822f
C114 net4 VPWR 1.16401f
C115 net6 _088_ 0.896031f
C116 _043_ _017_ 0.244201f
C117 a_8643_6249# VPWR 0.392083f
C118 net7 counter\[0\] 0.193184f
C119 _036_ _088_ 2.17834f
C120 _047_ _040_ 0.184738f
C121 net7 _008_ 0.551907f
C122 counter\[6\] net4 0.574581f
C123 counter\[5\] counter\[0\] 0.17228f
C124 counter\[6\] VPWR 2.11436f
C125 net1 _025_ 0.419365f
C126 a_2247_6575# VPWR 0.204902f
C127 counter\[10\] counter\[9\] 0.113039f
C128 net1 _092_ 0.211911f
C129 _090_ _030_ 0.491464f
C130 _059_ _080_ 0.16584f
C131 net3 clknet_0_clk 0.29246f
C132 a_6982_6005# VPWR 0.193556f
C133 a_8256_11177# _072_ 0.163988f
C134 counter\[0\] net9 0.46059f
C135 _026_ _073_ 0.779464f
C136 a_7791_9295# VPWR 0.191877f
C137 a_8643_6249# a_8779_6409# 0.136009f
C138 a_8779_6409# VPWR 0.17745f
C139 _086_ _068_ 0.121554f
C140 _049_ net13 0.190766f
C141 net9 _008_ 0.550319f
C142 _048_ net12 0.363638f
C143 a_7867_9019# VPWR 0.436471f
C144 _020_ net3 0.10769f
C145 a_6835_8751# clknet_1_1__leaf_clk 0.233938f
C146 a_4120_8731# _087_ 0.12321f
C147 _048_ _077_ 1.27586f
C148 net7 net10 0.17806f
C149 _043_ _053_ 0.119305f
C150 net5 _068_ 0.173676f
C151 net7 _084_ 0.104718f
C152 a_1731_6727# a_1827_6549# 0.310858f
C153 _005_ net1 0.233361f
C154 ready ones[7] 0.141229f
C155 a_6719_10615# VPWR 0.473656f
C156 a_8951_4949# VPWR 0.575618f
C157 a_8390_7119# clknet_1_1__leaf_clk 1.63485f
C158 _086_ _047_ 0.153868f
C159 _040_ a_4535_7232# 0.12488f
C160 _049_ _006_ 0.270876f
C161 net12 _022_ 0.107722f
C162 a_6425_10602# _045_ 0.222352f
C163 _015_ VPWR 2.38727f
C164 _069_ counter\[0\] 0.108299f
C165 _052_ net13 0.597326f
C166 _005_ net13 2.09319f
C167 _074_ _003_ 0.174401f
C168 _066_ _026_ 0.193441f
C169 _028_ _039_ 0.369055f
C170 _038_ counter\[1\] 0.186564f
C171 _039_ _091_ 0.151963f
C172 a_4307_8439# VPWR 0.210432f
C173 clknet_1_0__leaf_clk a_2118_6849# 0.455138f
C174 net1 _062_ 0.101961f
C175 net3 counter\[10\] 0.543441f
C176 clk _053_ 0.21925f
C177 counter\[4\] _000_ 0.403197f
C178 a_5142_3423# a_4535_3311# 0.136009f
C179 a_8999_5639# VPWR 0.388838f
C180 net9 _084_ 0.494968f
C181 _052_ _006_ 0.188052f
C182 counter\[3\] _073_ 0.1155f
C183 a_3847_8903# a_4120_8731# 0.167615f
C184 a_6375_6037# VPWR 0.447308f
C185 _016_ _046_ 0.188033f
C186 a_6423_11079# counter\[10\] 0.193426f
C187 a_1941_7125# _017_ 0.176818f
C188 _053_ _026_ 0.270508f
C189 a_8650_6153# _010_ 0.180854f
C190 net14 _087_ 0.527788f
C191 net5 counter\[7\] 0.384426f
C192 _069_ _084_ 1.18313f
C193 a_7442_8863# VPWR 0.179546f
C194 a_6375_6037# a_6982_6005# 0.136009f
C195 _034_ _021_ 0.80283f
C196 a_9091_10004# VPWR 0.278175f
C197 a_6361_3311# _003_ 0.114653f
C198 a_7189_8751# _022_ 0.114644f
C199 _070_ net13 0.641616f
C200 _037_ a_7663_7485# 0.192601f
C201 _068_ a_7111_4221# 0.164115f
C202 _023_ counter\[9\] 0.202106f
C203 _068_ a_1683_10496# 0.205089f
C204 clknet_0_clk a_8390_7119# 0.388577f
C205 a_6814_4765# VPWR 0.26014f
C206 a_10239_8751# net9 0.190764f
C207 _074_ _060_ 0.103692f
C208 _025_ _022_ 0.902837f
C209 a_7331_5853# a_6633_5487# 0.192261f
C210 a_1867_4399# _057_ 0.216013f
C211 a_5507_10357# VPWR 0.434986f
C212 clknet_1_0__leaf_clk counter\[3\] 0.280169f
C213 a_2866_3087# net8 0.182834f
C214 a_6987_2197# clknet_1_1__leaf_clk 0.221809f
C215 _090_ VPWR 0.646187f
C216 clknet_1_0__leaf_clk counter\[4\] 0.373806f
C217 net4 counter\[8\] 0.203989f
C218 net13 net8 0.372282f
C219 counter\[7\] clknet_1_1__leaf_clk 0.205951f
C220 net3 _035_ 1.43584f
C221 counter\[8\] VPWR 3.72486f
C222 _013_ _068_ 0.800684f
C223 _067_ counter\[1\] 1.05183f
C224 ones[9] ones[10] 0.178652f
C225 _002_ a_7725_10761# 0.121379f
C226 a_3799_10927# VPWR 0.234542f
C227 net9 _040_ 0.331992f
C228 a_4981_9991# VPWR 0.172207f
C229 _023_ net3 0.641295f
C230 net1 _088_ 0.245684f
C231 counter\[2\] _052_ 0.263272f
C232 _041_ _040_ 0.227694f
C233 _005_ counter\[2\] 0.417485f
C234 net6 _027_ 0.732173f
C235 net6 VPWR 2.35895f
C236 a_2313_4943# _018_ 0.115484f
C237 net14 net7 1.31451f
C238 net12 _024_ 0.216066f
C239 _039_ net4 0.109424f
C240 _036_ VPWR 0.633517f
C241 _066_ _001_ 1.18321f
C242 _033_ net8 0.692443f
C243 _039_ VPWR 1.86412f
C244 counter\[2\] _062_ 0.231496f
C245 net2 a_9096_4373# 0.204851f
C246 net3 counter\[1\] 0.311551f
C247 net7 net5 0.606654f
C248 _086_ counter\[5\] 0.102921f
C249 _034_ _033_ 0.240313f
C250 _085_ _042_ 0.130054f
C251 a_9586_6549# a_9515_6575# 0.239923f
C252 _063_ _047_ 0.101639f
C253 a_8631_2986# _008_ 0.109037f
C254 a_3413_2773# a_3854_2741# 0.110715f
C255 net5 counter\[5\] 0.350228f
C256 _077_ _073_ 0.111754f
C257 a_4234_2497# a_4227_2197# 0.962847f
C258 counter\[10\] _068_ 0.152807f
C259 net5 net9 1.37332f
C260 net1 _028_ 0.14089f
C261 a_9963_7663# ones[8] 0.112183f
C262 net5 _058_ 0.222477f
C263 a_8643_6249# a_8850_6308# 0.259379f
C264 net1 _091_ 0.520312f
C265 a_8850_6308# VPWR 0.245878f
C266 net5 _041_ 0.643791f
C267 _014_ net13 0.750341f
C268 a_9963_7663# VPWR 0.189628f
C269 _066_ net12 0.148661f
C270 _048_ net8 0.310045f
C271 a_4802_4132# VPWR 0.240829f
C272 _076_ net2 0.29981f
C273 a_9386_5761# _004_ 0.195142f
C274 counter\[2\] _031_ 0.178545f
C275 a_7407_6005# VPWR 0.416449f
C276 _002_ clknet_1_1__leaf_clk 0.149375f
C277 _072_ _073_ 0.729843f
C278 _054_ _082_ 0.131854f
C279 net7 clknet_1_1__leaf_clk 0.43514f
C280 _045_ _043_ 0.230894f
C281 a_8850_6308# a_8779_6409# 0.239923f
C282 a_8447_5175# _048_ 0.159275f
C283 a_4903_9295# _001_ 0.107548f
C284 a_9915_6337# VPWR 0.189423f
C285 _025_ _024_ 0.153001f
C286 _086_ _056_ 0.246598f
C287 a_7123_2223# a_6994_2497# 0.121264f
C288 _037_ net8 0.72111f
C289 net7 _093_ 0.288248f
C290 _028_ _033_ 0.259379f
C291 counter\[2\] net8 1.41362f
C292 _018_ net13 0.260473f
C293 _000_ _049_ 0.243521f
C294 clknet_1_0__leaf_clk net12 0.782915f
C295 a_1827_6549# a_2118_6849# 0.194892f
C296 clk net11 0.315547f
C297 a_5687_5175# _059_ 0.197894f
C298 _077_ _053_ 0.306169f
C299 a_7171_10601# VPWR 0.472489f
C300 a_8631_2986# _032_ 0.191109f
C301 a_6927_9301# counter\[0\] 0.423382f
C302 _061_ _092_ 0.237578f
C303 _037_ _034_ 0.137521f
C304 _058_ clknet_1_1__leaf_clk 0.24077f
C305 a_9595_3087# _039_ 0.105831f
C306 _021_ _027_ 0.157852f
C307 _093_ net9 0.970335f
C308 _021_ VPWR 0.834007f
C309 a_6633_5487# VPWR 0.292878f
C310 ready net9 0.15709f
C311 counter\[10\] _087_ 1.4542f
C312 _054_ VPWR 2.23804f
C313 _058_ _059_ 0.447438f
C314 _026_ net11 0.974094f
C315 _068_ _071_ 0.121638f
C316 counter\[6\] _021_ 0.361898f
C317 net1 _082_ 0.225085f
C318 a_9832_8181# VPWR 0.190828f
C319 counter\[0\] _060_ 0.69256f
C320 a_3697_6031# a_3797_6147# 0.167615f
C321 _076_ counter\[0\] 0.13891f
C322 a_6173_3311# _003_ 0.180545f
C323 _048_ _030_ 0.544073f
C324 net6 a_5507_10357# 0.136956f
C325 _069_ _093_ 0.984322f
C326 _071_ _047_ 0.674549f
C327 pulse rst 0.13211f
C328 ones[7] ones[2] 0.167004f
C329 counter\[9\] _038_ 0.119369f
C330 counter\[4\] _004_ 0.104057f
C331 _029_ counter\[0\] 0.10384f
C332 net7 clknet_0_clk 0.486405f
C333 _055_ _067_ 0.236563f
C334 _026_ _085_ 0.348682f
C335 _013_ a_6515_4074# 0.107904f
C336 a_7001_8751# a_6835_8751# 0.961627f
C337 ones[2] a_9871_2223# 0.109683f
C338 a_5675_4765# VPWR 0.187293f
C339 counter\[0\] _042_ 0.344661f
C340 a_3295_10615# a_3391_10615# 0.310858f
C341 _037_ _028_ 0.238149f
C342 clk rst 0.138937f
C343 a_6994_2497# VPWR 0.300469f
C344 net7 _020_ 0.820391f
C345 net1 VPWR 1.68089f
C346 counter\[2\] _028_ 0.119734f
C347 _068_ counter\[1\] 0.139356f
C348 counter\[4\] _074_ 0.14215f
C349 a_2866_3087# VPWR 0.214253f
C350 net6 _036_ 0.414566f
C351 net13 net4 0.495189f
C352 clknet_1_0__leaf_clk _049_ 0.107001f
C353 _043_ net2 0.13102f
C354 a_7239_4765# VPWR 0.179047f
C355 net13 VPWR 3.66744f
C356 _020_ counter\[5\] 0.551992f
C357 a_4073_7235# VPWR 0.211022f
C358 a_8175_6549# _053_ 0.138807f
C359 ones[8] _006_ 0.193744f
C360 a_5363_2880# VPWR 0.191126f
C361 counter\[1\] _047_ 0.244082f
C362 counter\[6\] net13 0.121344f
C363 a_4215_4087# VPWR 0.408137f
C364 net7 counter\[10\] 0.598152f
C365 a_6423_9991# a_6519_9813# 0.310858f
C366 a_9983_4917# a_9815_4943# 0.310858f
C367 _006_ VPWR 1.24918f
C368 _042_ net10 0.175405f
C369 _023_ counter\[7\] 0.337932f
C370 a_2382_7093# VPWR 0.190764f
C371 _084_ _042_ 1.3376f
C372 _033_ net4 0.644709f
C373 a_2555_10704# counter\[0\] 0.245586f
C374 net8 _024_ 0.253832f
C375 counter\[2\] _018_ 0.75771f
C376 net12 a_9687_7663# 0.184514f
C377 _033_ VPWR 1.72224f
C378 _026_ a_8720_8439# 0.137903f
C379 _023_ a_4535_7232# 0.168718f
C380 a_8256_11177# VPWR 0.169258f
C381 counter\[4\] _085_ 0.37483f
C382 _084_ ones[10] 0.154761f
C383 _089_ _060_ 0.331672f
C384 a_1460_9269# _059_ 0.182167f
C385 counter\[6\] _033_ 0.359715f
C386 net2 _026_ 0.11285f
C387 counter\[7\] counter\[1\] 0.276208f
C388 a_1775_7125# a_1941_7125# 0.966391f
C389 net3 a_10239_9839# 0.203175f
C390 _081_ VPWR 0.75228f
C391 _066_ _070_ 0.607665f
C392 _015_ net13 0.199169f
C393 a_1959_4949# _018_ 0.132481f
C394 _034_ _000_ 0.29901f
C395 ones[4] ones[0] 0.139374f
C396 _086_ _003_ 0.136682f
C397 ones[1] net8 0.193331f
C398 _087_ counter\[1\] 0.156104f
C399 _067_ counter\[9\] 0.231555f
C400 _066_ _031_ 0.473169f
C401 a_7419_5281# _087_ 0.115505f
C402 net12 a_6467_5487# 0.441289f
C403 a_2125_4949# a_2566_4917# 0.118966f
C404 _005_ a_3675_10601# 0.121026f
C405 a_3811_10761# a_3682_10505# 0.110715f
C406 _048_ _027_ 0.136893f
C407 _065_ counter\[0\] 0.195544f
C408 a_6810_10113# a_6939_9839# 0.119401f
C409 _048_ VPWR 1.09297f
C410 a_4227_2197# a_4434_2197# 0.273138f
C411 a_4234_2497# a_4363_2223# 0.110715f
C412 a_7307_10761# VPWR 0.198503f
C413 _044_ _026_ 0.27859f
C414 ones[5] _084_ 0.174409f
C415 _057_ VPWR 3.22826f
C416 counter\[3\] net2 1.34978f
C417 a_5141_4917# VPWR 0.197003f
C418 net3 counter\[9\] 0.226145f
C419 ones[6] _069_ 0.105121f
C420 _043_ net10 0.164471f
C421 a_4701_3311# VPWR 0.279655f
C422 _022_ VPWR 0.548234f
C423 _028_ _024_ 0.158066f
C424 _037_ VPWR 2.05219f
C425 _036_ _021_ 0.293467f
C426 counter\[0\] _026_ 0.134195f
C427 a_7039_3579# a_6871_3677# 0.310858f
C428 a_5717_4087# VPWR 0.15731f
C429 _064_ a_4903_9295# 0.185706f
C430 a_6927_9301# a_7534_9269# 0.136009f
C431 _074_ net12 0.310977f
C432 a_2318_6549# a_2111_6549# 0.273138f
C433 counter\[2\] VPWR 2.19658f
C434 net3 _067_ 0.455033f
C435 a_9435_9001# VPWR 0.489618f
C436 _040_ _042_ 0.270434f
C437 _053_ net8 0.201786f
C438 a_3611_4943# _060_ 0.259019f
C439 counter\[6\] _037_ 0.251734f
C440 counter\[5\] _035_ 1.28414f
C441 net9 _071_ 0.634122f
C442 net3 a_2971_8751# 0.102954f
C443 net12 net11 0.679168f
C444 a_6423_11079# counter\[9\] 0.237071f
C445 _019_ counter\[0\] 0.214875f
C446 net14 _060_ 0.437038f
C447 net14 _076_ 2.62277f
C448 a_7123_2223# a_7194_2197# 0.239923f
C449 _045_ _077_ 0.164652f
C450 _061_ _091_ 0.170694f
C451 a_4697_5461# clknet_0_clk 0.314925f
C452 _023_ counter\[5\] 0.822226f
C453 _028_ _073_ 0.401936f
C454 a_7407_4667# net3 0.16367f
C455 clknet_1_0__leaf_clk _034_ 0.552193f
C456 _043_ _032_ 1.25818f
C457 a_4602_3977# _020_ 0.370684f
C458 a_1959_4949# VPWR 0.463523f
C459 a_7001_8751# a_7699_9117# 0.192261f
C460 a_2118_6849# a_2111_6549# 0.962847f
C461 net7 counter\[1\] 0.150758f
C462 _070_ a_2603_10927# 0.196991f
C463 net5 _060_ 0.596416f
C464 _026_ net10 0.690381f
C465 ones[5] a_10239_8751# 0.116443f
C466 _023_ _041_ 0.116425f
C467 net1 a_4981_9991# 0.11457f
C468 net14 _042_ 0.380313f
C469 counter\[9\] _080_ 0.425929f
C470 a_6719_10615# counter\[2\] 0.128681f
C471 _055_ _068_ 2.20484f
C472 _093_ a_9096_4373# 0.123202f
C473 a_9386_5761# a_9379_5461# 0.965425f
C474 a_6906_5853# VPWR 0.268209f
C475 counter\[3\] counter\[0\] 0.563267f
C476 net1 net6 0.362812f
C477 counter\[2\] _015_ 0.383636f
C478 net2 _001_ 0.134654f
C479 _090_ _006_ 0.7767f
C480 counter\[4\] counter\[0\] 0.145399f
C481 _068_ _038_ 0.560514f
C482 a_6927_9301# clknet_1_1__leaf_clk 0.269581f
C483 _063_ a_3983_5056# 0.197084f
C484 _058_ counter\[1\] 0.774512f
C485 _067_ _080_ 0.131235f
C486 _086_ a_2460_3971# 0.10277f
C487 a_4771_2741# counter\[5\] 0.18874f
C488 a_4889_3311# _021_ 0.113517f
C489 a_6887_10615# a_7178_10505# 0.192261f
C490 counter\[0\] a_3431_4943# 0.243793f
C491 _043_ a_6169_6549# 0.213444f
C492 a_4123_9514# _089_ 0.197559f
C493 counter\[10\] _079_ 0.171889f
C494 clknet_1_0__leaf_clk _014_ 0.724666f
C495 _069_ counter\[1\] 0.112648f
C496 a_6375_4399# VPWR 0.449084f
C497 _039_ _006_ 1.02453f
C498 a_1867_4399# _074_ 0.115419f
C499 a_7274_9117# a_6835_8751# 0.260055f
C500 ones[2] net9 0.337653f
C501 net3 _080_ 0.359269f
C502 a_9197_6409# _010_ 0.114659f
C503 _009_ _047_ 0.386749f
C504 _055_ a_3247_2773# 0.442048f
C505 a_7194_2197# VPWR 0.24334f
C506 a_6283_7669# a_6475_7913# 0.101254f
C507 clk a_6169_6549# 0.306855f
C508 a_9503_8207# VPWR 0.241099f
C509 a_9815_4943# a_9117_4949# 0.194892f
C510 _029_ clknet_1_1__leaf_clk 0.135022f
C511 _059_ _060_ 0.726304f
C512 _067_ _050_ 2.29478f
C513 net6 _081_ 0.35043f
C514 a_4977_4399# VPWR 0.308114f
C515 net12 net2 0.111705f
C516 _024_ VPWR 1.45464f
C517 _042_ clknet_1_1__leaf_clk 0.593697f
C518 _005_ _045_ 0.342381f
C519 clknet_1_0__leaf_clk _018_ 0.139478f
C520 ones[7] net3 0.762288f
C521 _032_ counter\[3\] 0.691377f
C522 _000_ VPWR 0.560231f
C523 counter\[6\] _024_ 0.153509f
C524 counter\[7\] _011_ 0.122688f
C525 a_4595_4073# VPWR 0.401876f
C526 _086_ _043_ 0.409328f
C527 _057_ counter\[8\] 0.110781f
C528 a_2807_7093# VPWR 0.416761f
C529 _061_ VPWR 0.304653f
C530 ones[8] ones[1] 0.205179f
C531 counter\[9\] _068_ 0.413676f
C532 _013_ a_4234_2497# 0.18425f
C533 a_6871_3677# VPWR 0.212701f
C534 _073_ VPWR 1.85528f
C535 _090_ counter\[2\] 0.350035f
C536 _037_ counter\[8\] 1.53321f
C537 _006_ a_7541_2223# 0.119626f
C538 _090_ a_9435_9001# 0.191107f
C539 a_5717_4087# counter\[8\] 0.178306f
C540 a_1670_6351# _049_ 0.150691f
C541 ones[1] VPWR 0.138934f
C542 counter\[2\] counter\[8\] 0.738451f
C543 net6 _057_ 0.131928f
C544 a_8447_8916# VPWR 0.212977f
C545 _044_ net12 1.06468f
C546 counter\[9\] _047_ 0.683142f
C547 _017_ VPWR 0.411041f
C548 _074_ _070_ 0.129746f
C549 net14 _026_ 0.603968f
C550 _021_ net13 0.16434f
C551 _063_ _060_ 0.323923f
C552 _066_ VPWR 0.967442f
C553 _054_ net13 0.41802f
C554 a_4595_4073# _015_ 0.442035f
C555 counter\[2\] _039_ 0.285377f
C556 _029_ clknet_0_clk 0.50049f
C557 a_2566_4917# a_2398_4943# 0.239923f
C558 net3 _068_ 0.10018f
C559 _025_ net2 0.104581f
C560 net2 _049_ 0.243096f
C561 a_7010_9813# a_6939_9839# 0.239923f
C562 _054_ _006_ 0.301181f
C563 _055_ net7 0.281559f
C564 a_3123_6031# VPWR 0.201102f
C565 _043_ clknet_1_1__leaf_clk 0.144978f
C566 a_4434_2197# a_4363_2223# 0.239923f
C567 _074_ net8 0.12717f
C568 ones[0] a_10239_9839# 0.108562f
C569 _079_ counter\[1\] 0.260103f
C570 _053_ VPWR 0.898184f
C571 clknet_1_0__leaf_clk VPWR 5.62373f
C572 net5 _019_ 0.150716f
C573 _070_ _085_ 0.227067f
C574 ready pulse 0.129624f
C575 counter\[10\] _060_ 0.1304f
C576 a_6814_4765# a_6375_4399# 0.260055f
C577 a_6982_4511# a_6541_4399# 0.119401f
C578 a_9079_3855# a_9247_3829# 0.310858f
C579 a_10239_10927# VPWR 0.275085f
C580 a_2991_4917# a_2823_4943# 0.310858f
C581 a_1461_9813# net12 0.171646f
C582 a_4974_3677# VPWR 0.24224f
C583 counter\[6\] _053_ 0.168276f
C584 clknet_1_0__leaf_clk counter\[6\] 0.382918f
C585 a_6541_6037# _001_ 0.226837f
C586 _074_ _034_ 0.198027f
C587 _065_ clknet_1_1__leaf_clk 0.12542f
C588 clk clknet_1_1__leaf_clk 1.57728f
C589 _021_ _081_ 0.626704f
C590 net14 counter\[3\] 0.167681f
C591 a_9386_5761# clknet_1_1__leaf_clk 0.422786f
C592 a_8381_3861# a_8822_3829# 0.114265f
C593 a_8459_4551# VPWR 0.213124f
C594 _045_ _034_ 0.212834f
C595 counter\[5\] _011_ 0.331496f
C596 _062_ net2 0.255637f
C597 _088_ net11 0.138263f
C598 a_7847_3855# net11 0.190109f
C599 _086_ counter\[4\] 0.145486f
C600 a_6810_10113# a_6803_9813# 0.961981f
C601 a_4111_2767# a_3413_2773# 0.189491f
C602 net5 counter\[3\] 0.363251f
C603 a_3431_4943# a_3611_4943# 0.185422f
C604 ones[3] a_10239_7663# 0.110226f
C605 _026_ clknet_1_1__leaf_clk 0.151216f
C606 a_7171_10601# a_7307_10761# 0.136009f
C607 _068_ _080_ 0.108916f
C608 a_6994_2497# _006_ 0.181793f
C609 net5 counter\[4\] 0.275844f
C610 a_4903_9295# VPWR 0.255617f
C611 net12 _032_ 0.287211f
C612 a_4215_4087# net13 0.107867f
C613 net1 _033_ 0.245874f
C614 _014_ a_3413_2773# 0.562455f
C615 _058_ a_9739_6005# 0.189565f
C616 _019_ clknet_1_1__leaf_clk 0.195945f
C617 a_3675_10601# VPWR 0.705368f
C618 _033_ net13 0.205735f
C619 a_2603_10927# VPWR 0.238855f
C620 a_9386_5761# a_9515_5487# 0.110715f
C621 a_9379_5461# a_9586_5461# 0.273138f
C622 _055_ _056_ 0.11855f
C623 a_10147_4399# VPWR 0.196408f
C624 _043_ clknet_0_clk 0.492309f
C625 a_4701_3311# _021_ 0.18054f
C626 a_7663_7485# net10 0.154259f
C627 a_9305_4943# _016_ 0.114807f
C628 _074_ _028_ 0.203327f
C629 a_2509_4663# VPWR 0.200625f
C630 a_6173_3311# a_6614_3423# 0.110715f
C631 a_9379_6549# a_9515_6575# 0.141453f
C632 a_9386_6849# _007_ 0.180673f
C633 _071_ _060_ 1.07238f
C634 _014_ net11 0.124166f
C635 _028_ net11 0.218777f
C636 a_7093_9301# a_7534_9269# 0.110715f
C637 _025_ net10 0.334553f
C638 net5 a_7093_9301# 0.422395f
C639 net2 _031_ 0.1045f
C640 _073_ counter\[8\] 0.615244f
C641 _007_ clknet_1_1__leaf_clk 0.182923f
C642 _077_ a_4668_7913# 0.106122f
C643 a_2787_8207# VPWR 0.262992f
C644 a_9832_8181# counter\[2\] 0.145695f
C645 _049_ _084_ 0.116904f
C646 counter\[0\] _062_ 0.171585f
C647 counter\[5\] counter\[9\] 0.391834f
C648 ones[8] a_9687_7663# 0.110357f
C649 net7 _067_ 0.231354f
C650 net6 _061_ 0.346693f
C651 _044_ _064_ 0.123095f
C652 _062_ _008_ 0.694383f
C653 net5 _001_ 0.443975f
C654 net12 _040_ 0.106546f
C655 _023_ _060_ 0.116757f
C656 a_10239_10383# ones[4] 0.110639f
C657 a_5359_4943# counter\[4\] 0.103687f
C658 counter\[4\] _093_ 1.1902f
C659 a_1499_5056# _068_ 0.203093f
C660 a_3682_10505# counter\[1\] 0.264209f
C661 _058_ counter\[9\] 0.257308f
C662 a_9687_7663# VPWR 0.252119f
C663 net7 _078_ 0.518435f
C664 _026_ clknet_0_clk 0.116344f
C665 _066_ _090_ 0.103941f
C666 _039_ _073_ 0.227449f
C667 _014_ _085_ 0.453584f
C668 counter\[9\] _041_ 0.139942f
C669 ones[4] ones[10] 0.1711f
C670 a_7939_6031# net10 0.18966f
C671 net1 _022_ 0.558673f
C672 a_6541_4399# _011_ 0.183699f
C673 _034_ net2 0.368583f
C674 _028_ a_9687_4399# 0.169219f
C675 a_5250_4765# VPWR 0.250391f
C676 net1 _037_ 0.151947f
C677 net3 _002_ 0.4481f
C678 net7 net3 0.327318f
C679 net1 counter\[2\] 0.232621f
C680 clk counter\[10\] 0.324012f
C681 _069_ counter\[9\] 0.186198f
C682 _062_ _084_ 0.117366f
C683 ones[6] _043_ 0.196902f
C684 counter\[5\] net3 1.13362f
C685 _029_ counter\[1\] 0.138388f
C686 counter\[2\] net13 0.367914f
C687 a_5785_9813# VPWR 0.232058f
C688 a_9390_4943# VPWR 0.252873f
C689 a_6835_8751# _087_ 0.426305f
C690 counter\[0\] _031_ 0.775454f
C691 a_6467_5487# VPWR 0.483307f
C692 counter\[1\] _042_ 0.514354f
C693 a_4595_4073# a_4802_4132# 0.260055f
C694 counter\[9\] _056_ 0.839614f
C695 a_9213_3463# VPWR 0.164909f
C696 _058_ net3 0.543699f
C697 a_9225_4649# VPWR 0.189894f
C698 net5 net12 0.410238f
C699 counter\[2\] _006_ 0.448644f
C700 _037_ _033_ 0.101372f
C701 a_9435_9001# _006_ 0.112318f
C702 _019_ a_6007_8207# 0.108698f
C703 a_2879_3855# _088_ 0.129023f
C704 a_3697_6031# _080_ 0.150764f
C705 _044_ _034_ 0.181206f
C706 counter\[2\] _033_ 0.187702f
C707 _004_ VPWR 0.489613f
C708 counter\[4\] clknet_0_clk 0.517612f
C709 a_3413_2773# VPWR 0.302469f
C710 a_9079_3855# VPWR 0.176721f
C711 a_9963_7663# ones[1] 0.110384f
C712 net2 _030_ 0.12162f
C713 _020_ counter\[3\] 0.333787f
C714 a_9095_6549# a_9386_6849# 0.194623f
C715 _014_ net2 0.293586f
C716 ones[9] VPWR 0.383591f
C717 _083_ VPWR 0.488251f
C718 _028_ net2 0.696159f
C719 a_8907_2986# VPWR 0.223476f
C720 counter\[4\] _020_ 0.112351f
C721 a_9390_4943# a_8951_4949# 0.273138f
C722 _074_ VPWR 3.5737f
C723 _018_ a_2125_4949# 0.261658f
C724 net11 net4 0.259135f
C725 counter\[5\] _080_ 0.136816f
C726 net11 VPWR 1.27521f
C727 a_1867_3561# VPWR 0.241733f
C728 a_1827_6549# VPWR 0.213595f
C729 _074_ counter\[6\] 0.790133f
C730 _045_ VPWR 2.53168f
C731 a_8447_8439# a_8720_8439# 0.167615f
C732 a_8569_3855# _015_ 0.114816f
C733 net12 clknet_1_1__leaf_clk 0.280938f
C734 ones[7] net7 0.122798f
C735 net14 _025_ 0.261897f
C736 net14 _092_ 0.137123f
C737 _087_ _047_ 0.227829f
C738 net12 _093_ 0.381929f
C739 net7 a_10239_7663# 0.208504f
C740 a_6803_9813# clknet_1_1__leaf_clk 0.290418f
C741 _086_ _049_ 2.80824f
C742 _044_ _028_ 0.192321f
C743 a_5675_4765# a_4977_4399# 0.194892f
C744 _026_ _071_ 0.195764f
C745 net7 a_8390_7119# 0.285011f
C746 _085_ VPWR 0.539997f
C747 net5 _025_ 0.328599f
C748 _020_ a_10195_7338# 0.107531f
C749 a_8822_3829# a_8654_3855# 0.239923f
C750 a_9687_4399# VPWR 0.185194f
C751 _028_ counter\[0\] 0.739841f
C752 _015_ net11 0.188529f
C753 _064_ _040_ 0.67874f
C754 a_6803_9813# a_7010_9813# 0.260055f
C755 a_5399_3677# a_5567_3579# 0.310858f
C756 _065_ counter\[1\] 0.115863f
C757 a_7178_10505# _002_ 0.243147f
C758 net2 _082_ 0.103746f
C759 a_9961_8207# VPWR 0.204065f
C760 a_1670_6351# VPWR 0.201113f
C761 _005_ net5 0.103677f
C762 ones[10] a_9687_10927# 0.120688f
C763 net14 _062_ 0.284973f
C764 a_1775_7125# VPWR 0.744008f
C765 a_1499_5056# counter\[5\] 0.238679f
C766 rst VPWR 0.19347f
C767 a_3882_10660# VPWR 0.245645f
C768 a_9515_6575# VPWR 0.181951f
C769 a_2125_4949# VPWR 0.314919f
C770 _021_ _053_ 0.397234f
C771 clknet_1_0__leaf_clk _021_ 0.269379f
C772 net7 _068_ 0.128855f
C773 _026_ counter\[1\] 0.104559f
C774 a_9586_5461# a_9515_5487# 0.239923f
C775 a_3601_2767# _014_ 0.124776f
C776 a_4227_2197# VPWR 0.615265f
C777 a_8720_8439# VPWR 0.164599f
C778 counter\[9\] a_1731_6727# 0.124437f
C779 _055_ _060_ 0.310604f
C780 counter\[4\] _071_ 0.228663f
C781 _023_ a_3029_6031# 0.121122f
C782 counter\[5\] _068_ 0.223659f
C783 _091_ _084_ 0.147855f
C784 ones[3] _069_ 0.14545f
C785 _063_ net12 0.439882f
C786 a_4227_2197# counter\[6\] 0.148982f
C787 a_6614_3423# a_6446_3677# 0.239923f
C788 net2 VPWR 3.30604f
C789 _020_ net12 0.172566f
C790 a_6927_9301# _012_ 0.120808f
C791 a_6729_4399# _011_ 0.113498f
C792 net5 _064_ 0.113399f
C793 _044_ _082_ 0.80509f
C794 a_2823_4943# VPWR 0.199433f
C795 a_4521_8903# _025_ 0.123607f
C796 ones[1] _006_ 0.114005f
C797 _006_ a_8447_8916# 0.133636f
C798 _032_ _030_ 0.170317f
C799 _029_ _038_ 0.624335f
C800 _005_ clknet_1_1__leaf_clk 0.120039f
C801 _034_ _040_ 0.1008f
C802 _066_ a_5363_2880# 0.194827f
C803 _061_ _081_ 0.419111f
C804 _067_ _003_ 0.394661f
C805 counter\[3\] counter\[1\] 1.06295f
C806 a_9933_6575# _007_ 0.113637f
C807 net1 _053_ 0.497475f
C808 a_2879_3855# VPWR 0.211165f
C809 counter\[4\] counter\[1\] 0.225836f
C810 a_4697_5461# _080_ 0.191915f
C811 _039_ _004_ 0.135732f
C812 clknet_1_0__leaf_clk net13 0.206219f
C813 counter\[5\] counter\[7\] 0.338288f
C814 _057_ _024_ 0.145607f
C815 _044_ VPWR 1.00911f
C816 net7 a_7847_3133# 0.223983f
C817 a_10239_10927# net13 0.21399f
C818 _069_ _047_ 0.628907f
C819 a_7366_9295# a_7534_9269# 0.239923f
C820 net5 net8 0.201742f
C821 net14 _034_ 0.218483f
C822 _037_ _024_ 0.241533f
C823 _058_ counter\[7\] 0.665026f
C824 counter\[0\] net4 0.144987f
C825 a_6519_9813# VPWR 0.194163f
C826 a_9815_4943# VPWR 0.185763f
C827 counter\[0\] VPWR 5.18572f
C828 a_4771_2741# counter\[4\] 0.159501f
C829 net6 net11 0.142364f
C830 a_2787_8207# _021_ 0.101844f
C831 _008_ net4 0.188184f
C832 _033_ _053_ 0.556375f
C833 _008_ VPWR 0.920542f
C834 _063_ _049_ 1.00229f
C835 a_4602_3977# a_4731_4233# 0.118966f
C836 _039_ net11 0.223222f
C837 _064_ _059_ 1.73876f
C838 _045_ _036_ 0.375551f
C839 _028_ _040_ 0.31527f
C840 _020_ _092_ 0.448845f
C841 a_8215_10496# _031_ 0.220248f
C842 a_2879_3855# _015_ 0.10736f
C843 _031_ clknet_1_1__leaf_clk 0.336217f
C844 a_9386_6849# a_9379_6549# 0.966678f
C845 a_1461_9813# VPWR 0.214667f
C846 _069_ _087_ 0.185879f
C847 net10 VPWR 4.00797f
C848 counter\[9\] _042_ 0.625199f
C849 _084_ VPWR 1.57132f
C850 a_9379_6549# clknet_1_1__leaf_clk 0.303855f
C851 a_8381_3861# VPWR 0.279675f
C852 counter\[0\] _015_ 0.283706f
C853 _003_ _080_ 0.179957f
C854 a_6810_10113# VPWR 0.294428f
C855 net14 _014_ 0.367858f
C856 _063_ _062_ 0.285806f
C857 net14 _028_ 0.267183f
C858 a_4535_3311# VPWR 0.447487f
C859 net14 _091_ 0.242669f
C860 a_2111_6549# VPWR 0.653635f
C861 a_6703_2197# a_6607_2375# 0.310858f
C862 a_2460_3971# counter\[9\] 0.196461f
C863 _043_ _009_ 0.155235f
C864 net3 _060_ 0.259995f
C865 clk _038_ 0.187921f
C866 _023_ net12 0.174136f
C867 a_6467_5487# a_6633_5487# 0.963608f
C868 a_9379_5461# VPWR 0.673727f
C869 a_2247_6575# a_2111_6549# 0.141453f
C870 _005_ counter\[10\] 0.126236f
C871 _032_ net4 0.453024f
C872 a_6173_3311# VPWR 0.297552f
C873 net7 counter\[5\] 0.138369f
C874 _046_ net12 0.679344f
C875 _032_ VPWR 0.839959f
C876 _029_ net3 0.189488f
C877 clknet_1_0__leaf_clk a_4701_3311# 0.483374f
C878 _016_ _043_ 0.90032f
C879 a_10195_7338# _051_ 0.191227f
C880 _009_ a_2118_6849# 0.183713f
C881 _089_ VPWR 0.489449f
C882 net7 net9 1.20276f
C883 _038_ _026_ 0.110278f
C884 net3 _042_ 0.375291f
C885 net12 counter\[1\] 0.840744f
C886 net7 a_7980_4649# 0.166029f
C887 _076_ _075_ 0.571351f
C888 _086_ _018_ 0.125631f
C889 a_8822_3829# a_8215_3861# 0.136001f
C890 a_8381_3861# _015_ 0.255024f
C891 a_10239_8751# VPWR 0.213289f
C892 a_6541_6037# VPWR 0.284751f
C893 a_4811_4399# a_5418_4511# 0.141453f
C894 _058_ counter\[5\] 0.579854f
C895 ones[6] a_7939_6031# 0.108611f
C896 _019_ _038_ 0.88903f
C897 a_4123_9514# _009_ 0.109575f
C898 a_4120_8731# VPWR 0.174101f
C899 clknet_1_0__leaf_clk a_1959_4949# 0.216845f
C900 _028_ a_8215_10496# 0.176292f
C901 _030_ clknet_1_1__leaf_clk 0.639301f
C902 a_4977_4399# _000_ 0.180554f
C903 a_4668_7913# VPWR 0.16471f
C904 a_6541_6037# a_6982_6005# 0.124191f
C905 _028_ clknet_1_1__leaf_clk 0.257839f
C906 a_6169_6549# VPWR 1.26082f
C907 counter\[6\] a_4668_7913# 0.169431f
C908 a_9503_8207# _073_ 0.18599f
C909 a_9386_5761# a_9095_5461# 0.194892f
C910 a_2398_4943# VPWR 0.255099f
C911 _040_ VPWR 1.03067f
C912 _020_ net8 1.9209f
C913 a_4311_4087# a_4602_3977# 0.192261f
C914 a_4363_2223# VPWR 0.182281f
C915 a_3811_10761# VPWR 0.177734f
C916 a_2879_3855# _036_ 0.196751f
C917 counter\[6\] _040_ 0.190423f
C918 counter\[10\] _031_ 0.173326f
C919 counter\[4\] _038_ 0.152198f
C920 _042_ _080_ 0.102024f
C921 a_7239_6031# VPWR 0.17932f
C922 a_4627_5056# _060_ 0.175363f
C923 counter\[0\] counter\[8\] 0.624978f
C924 counter\[3\] _011_ 0.151747f
C925 a_4279_2741# a_4111_2767# 0.310858f
C926 a_3611_4943# VPWR 0.168658f
C927 counter\[4\] _011_ 0.25068f
C928 _058_ _056_ 0.107591f
C929 _006_ _004_ 0.132511f
C930 _043_ net3 0.140647f
C931 _074_ net13 0.121901f
C932 net14 VPWR 1.83646f
C933 clknet_1_0__leaf_clk a_6375_4399# 0.214763f
C934 net1 _045_ 0.886487f
C935 a_2682_3311# counter\[7\] 0.170585f
C936 counter\[0\] _039_ 0.378719f
C937 clk _078_ 0.21372f
C938 _086_ VPWR 1.97318f
C939 a_6375_6037# a_6541_6037# 0.966899f
C940 a_7290_7119# VPWR 0.214734f
C941 a_9915_6337# net2 0.211132f
C942 net5 _027_ 0.141624f
C943 _090_ _084_ 0.226844f
C944 a_6007_3311# counter\[3\] 0.328063f
C945 a_7534_9269# VPWR 0.182212f
C946 _045_ a_4073_7235# 0.12997f
C947 net5 VPWR 3.93133f
C948 a_2971_8751# _026_ 0.113463f
C949 _084_ counter\[8\] 0.116885f
C950 clknet_1_0__leaf_clk a_4977_4399# 0.460216f
C951 counter\[7\] _003_ 0.106066f
C952 a_8393_6825# VPWR 0.281951f
C953 net5 counter\[6\] 0.476233f
C954 _053_ _024_ 0.204634f
C955 _082_ clknet_1_1__leaf_clk 0.413226f
C956 net14 a_7867_9019# 0.202296f
C957 a_4234_2497# _068_ 0.454649f
C958 _033_ net11 0.143455f
C959 net6 net10 0.196441f
C960 _063_ _091_ 0.535163f
C961 clknet_1_0__leaf_clk _000_ 0.504266f
C962 _062_ counter\[1\] 0.122246f
C963 clknet_1_0__leaf_clk a_4595_4073# 0.308384f
C964 _020_ _028_ 0.151829f
C965 net3 _026_ 0.697403f
C966 counter\[3\] counter\[9\] 0.142698f
C967 _020_ _091_ 0.240464f
C968 _090_ _032_ 0.281828f
C969 _074_ _081_ 0.568052f
C970 _054_ net2 0.564281f
C971 a_6283_7669# _031_ 0.128487f
C972 _043_ _080_ 0.471965f
C973 _012_ a_7093_9301# 0.269864f
C974 counter\[4\] counter\[9\] 0.665946f
C975 _005_ ones[2] 0.818225f
C976 counter\[2\] a_5785_9813# 0.20178f
C977 _060_ _047_ 1.00462f
C978 a_9386_6849# VPWR 0.305921f
C979 _016_ a_9117_4949# 0.25859f
C980 a_8215_10496# VPWR 0.202662f
C981 a_3847_2375# a_3943_2197# 0.310858f
C982 a_8643_6249# clknet_1_1__leaf_clk 0.731607f
C983 a_1670_6351# net13 0.180018f
C984 counter\[4\] _067_ 0.196983f
C985 counter\[10\] _028_ 1.04513f
C986 clknet_1_1__leaf_clk VPWR 6.18245f
C987 a_7886_3311# net9 0.121002f
C988 counter\[3\] _078_ 0.307649f
C989 _035_ net8 0.803972f
C990 _055_ net12 1.56929f
C991 a_5359_4943# VPWR 0.202857f
C992 _093_ VPWR 1.30536f
C993 ready VPWR 0.209082f
C994 _078_ a_9091_8439# 0.195814f
C995 _047_ _042_ 0.134962f
C996 _059_ VPWR 0.902677f
C997 _074_ _057_ 0.122958f
C998 a_7111_4221# VPWR 0.459362f
C999 _023_ net8 0.859238f
C1000 a_4521_8903# VPWR 0.145584f
C1001 a_8654_3855# VPWR 0.253036f
C1002 net3 counter\[3\] 0.763275f
C1003 a_1683_10496# VPWR 0.267205f
C1004 ones[3] ones[5] 0.172207f
C1005 a_1775_7125# a_2382_7093# 0.141453f
C1006 a_3295_10615# VPWR 0.427721f
C1007 counter\[7\] _060_ 0.623997f
C1008 _083_ a_5717_4087# 0.10615f
C1009 net1 net2 0.294402f
C1010 a_7010_9813# VPWR 0.257172f
C1011 counter\[4\] net3 0.112988f
C1012 _074_ _037_ 1.04855f
C1013 counter\[10\] _018_ 0.282343f
C1014 net12 _011_ 0.112718f
C1015 a_7407_6005# net10 0.118905f
C1016 counter\[0\] _021_ 0.128714f
C1017 ones[7] clk 0.245378f
C1018 _023_ _034_ 0.363644f
C1019 _087_ _060_ 0.202746f
C1020 _045_ _022_ 0.394338f
C1021 a_6467_5487# a_6906_5853# 0.260055f
C1022 a_9515_5487# VPWR 0.180125f
C1023 a_8951_4949# clknet_1_1__leaf_clk 0.225991f
C1024 counter\[2\] net11 0.242369f
C1025 a_6446_3677# VPWR 0.248799f
C1026 _045_ counter\[2\] 0.330314f
C1027 a_4279_2741# VPWR 0.395685f
C1028 net2 _006_ 0.372787f
C1029 net6 _040_ 0.461107f
C1030 counter\[4\] _075_ 0.733532f
C1031 _013_ VPWR 0.546809f
C1032 _033_ net2 0.191969f
C1033 a_3029_6031# _080_ 0.109365f
C1034 a_7847_3133# _042_ 0.111643f
C1035 _013_ counter\[6\] 0.404548f
C1036 clknet_0_clk net4 0.178041f
C1037 _037_ _085_ 0.917964f
C1038 a_2191_10615# counter\[1\] 0.182977f
C1039 clknet_0_clk VPWR 2.44763f
C1040 a_10199_2197# VPWR 0.355224f
C1041 a_3797_6147# VPWR 0.204009f
C1042 _020_ ones[8] 0.151118f
C1043 _063_ net4 0.843224f
C1044 a_6375_6037# clknet_1_1__leaf_clk 0.734594f
C1045 _063_ VPWR 0.595405f
C1046 a_3847_8903# _060_ 0.131175f
C1047 _086_ counter\[8\] 0.116134f
C1048 _044_ a_4073_7235# 0.212542f
C1049 net14 a_4981_9991# 0.163162f
C1050 a_6994_2497# counter\[0\] 0.328982f
C1051 net1 counter\[0\] 0.140463f
C1052 _020_ VPWR 0.894029f
C1053 a_3847_2375# VPWR 0.399067f
C1054 _055_ a_1867_4399# 0.165196f
C1055 _065_ _068_ 0.241547f
C1056 _023_ _028_ 0.209849f
C1057 net12 counter\[9\] 0.134418f
C1058 net14 _039_ 0.138086f
C1059 a_6614_3423# a_6007_3311# 0.136009f
C1060 clknet_1_0__leaf_clk a_3675_10601# 0.236089f
C1061 ones[6] _082_ 0.32864f
C1062 _046_ _028_ 0.126863f
C1063 a_6007_8207# VPWR 0.260799f
C1064 _055_ _052_ 0.176658f
C1065 _011_ _092_ 0.693892f
C1066 net6 net5 0.646643f
C1067 a_9503_8207# _004_ 0.111666f
C1068 net5 _036_ 0.762591f
C1069 counter\[10\] VPWR 1.97082f
C1070 net7 _060_ 0.156624f
C1071 a_3854_2741# a_3247_2773# 0.136009f
C1072 net5 _039_ 0.564399f
C1073 counter\[0\] _006_ 0.358419f
C1074 _028_ counter\[1\] 0.154408f
C1075 _068_ _026_ 0.132055f
C1076 a_8263_6263# VPWR 0.38207f
C1077 _091_ counter\[1\] 0.136294f
C1078 _033_ counter\[0\] 1.79157f
C1079 _006_ _008_ 0.406029f
C1080 net1 net10 0.336355f
C1081 _043_ counter\[7\] 0.350362f
C1082 counter\[5\] _060_ 0.453407f
C1083 _025_ _012_ 0.705139f
C1084 net1 _084_ 0.374645f
C1085 ones[6] ones[8] 0.231126f
C1086 _078_ _077_ 0.133365f
C1087 a_10287_6250# _007_ 0.13499f
C1088 _026_ _047_ 0.241799f
C1089 counter\[9\] _072_ 0.590795f
C1090 _038_ _062_ 0.198861f
C1091 a_7407_6005# a_7239_6031# 0.310858f
C1092 _084_ net13 2.43573f
C1093 _076_ net9 0.131921f
C1094 net7 _042_ 0.11269f
C1095 _058_ _060_ 0.456995f
C1096 ones[6] VPWR 0.188981f
C1097 a_6987_2197# _065_ 0.508766f
C1098 counter\[0\] _081_ 0.127363f
C1099 a_1959_4949# a_2125_4949# 0.965735f
C1100 _074_ _024_ 0.48218f
C1101 a_4595_4073# _083_ 0.106912f
C1102 _029_ a_6515_4074# 0.187311f
C1103 counter\[5\] _042_ 0.133077f
C1104 a_1499_5056# counter\[4\] 0.105725f
C1105 _066_ a_5785_9813# 0.114542f
C1106 net3 a_6803_9813# 0.470962f
C1107 a_3391_10615# a_3682_10505# 0.192122f
C1108 a_6391_2767# _028_ 0.191907f
C1109 clk _087_ 0.14308f
C1110 a_1683_10496# counter\[8\] 0.217664f
C1111 counter\[3\] _068_ 2.85303f
C1112 _039_ clknet_1_1__leaf_clk 0.78272f
C1113 net5 a_9963_7663# 0.199466f
C1114 ones[0] ones[5] 0.120241f
C1115 counter\[9\] _049_ 0.141384f
C1116 counter\[4\] _068_ 0.747871f
C1117 _016_ _062_ 0.127926f
C1118 _048_ counter\[0\] 0.127749f
C1119 _093_ _039_ 0.358359f
C1120 a_8359_6263# VPWR 0.181073f
C1121 _071_ _027_ 0.328415f
C1122 net1 a_6541_6037# 0.107855f
C1123 ones[4] VPWR 0.441833f
C1124 a_7847_3133# _026_ 0.145534f
C1125 counter\[3\] _047_ 0.155877f
C1126 _071_ VPWR 0.918728f
C1127 clknet_1_0__leaf_clk a_6467_5487# 0.221971f
C1128 _082_ counter\[1\] 0.339297f
C1129 counter\[6\] _071_ 0.124751f
C1130 net12 _080_ 0.130789f
C1131 _037_ counter\[0\] 0.461197f
C1132 _035_ VPWR 1.60396f
C1133 counter\[2\] counter\[0\] 0.427445f
C1134 a_7959_9269# VPWR 0.410379f
C1135 net1 a_6169_6549# 0.115864f
C1136 _023_ VPWR 1.62968f
C1137 counter\[2\] _008_ 1.4534f
C1138 _067_ _052_ 0.922451f
C1139 _066_ _045_ 0.159223f
C1140 counter\[9\] _062_ 0.175916f
C1141 net7 _043_ 0.39625f
C1142 net3 _049_ 0.465358f
C1143 _046_ VPWR 0.700186f
C1144 clknet_1_0__leaf_clk _083_ 0.456727f
C1145 a_6375_4399# net2 0.428991f
C1146 ones[9] a_10239_10927# 0.110649f
C1147 counter\[4\] counter\[7\] 0.922486f
C1148 counter\[1\] net4 1.51825f
C1149 a_7959_9269# a_7791_9295# 0.310858f
C1150 a_8215_3861# VPWR 0.59979f
C1151 clknet_1_0__leaf_clk _074_ 1.44088f
C1152 _022_ net10 0.239795f
C1153 a_1460_9269# _060_ 0.1787f
C1154 counter\[1\] VPWR 2.63774f
C1155 _010_ _082_ 0.267909f
C1156 _037_ net10 0.901434f
C1157 a_7419_5281# VPWR 0.213379f
C1158 net7 _065_ 0.400344f
C1159 net7 clk 0.159393f
C1160 _039_ clknet_0_clk 0.343934f
C1161 clknet_1_0__leaf_clk net11 0.324747f
C1162 _043_ net9 0.181355f
C1163 _066_ _085_ 0.215064f
C1164 _050_ net12 0.408913f
C1165 _058_ _043_ 0.117401f
C1166 _043_ _041_ 0.528713f
C1167 a_8381_3861# counter\[2\] 0.265296f
C1168 a_4701_3311# a_4535_3311# 0.961627f
C1169 a_8109_5639# VPWR 0.166439f
C1170 a_9435_9001# _084_ 0.102421f
C1171 _063_ _039_ 0.39856f
C1172 a_1501_6031# VPWR 0.234447f
C1173 net6 a_3847_2375# 0.102786f
C1174 _048_ _032_ 1.34738f
C1175 counter\[2\] a_6810_10113# 0.10118f
C1176 net14 net1 1.1063f
C1177 _090_ counter\[10\] 0.361387f
C1178 a_7171_10601# clknet_1_1__leaf_clk 0.296424f
C1179 counter\[10\] counter\[8\] 0.232798f
C1180 a_4627_6031# VPWR 0.194759f
C1181 ones[8] _010_ 0.390012f
C1182 net7 _026_ 1.45172f
C1183 a_8459_4551# net11 0.120474f
C1184 a_4771_2741# VPWR 0.395132f
C1185 ones[2] VPWR 0.734082f
C1186 _086_ net13 0.363375f
C1187 _067_ _070_ 0.149016f
C1188 a_3187_2251# _080_ 0.111987f
C1189 a_4771_2741# counter\[6\] 0.122377f
C1190 _054_ clknet_1_1__leaf_clk 0.345065f
C1191 _010_ VPWR 0.433874f
C1192 _049_ _080_ 0.177776f
C1193 a_6391_2767# VPWR 0.441771f
C1194 a_7001_8751# VPWR 0.311468f
C1195 a_8215_3861# _015_ 0.112695f
C1196 net14 _006_ 0.104826f
C1197 counter\[10\] _039_ 0.191619f
C1198 net3 _064_ 0.344885f
C1199 _028_ _038_ 0.114656f
C1200 net14 _033_ 0.12762f
C1201 _026_ a_7980_4649# 0.100729f
C1202 _062_ _075_ 0.301437f
C1203 _051_ VPWR 0.579975f
C1204 clk _069_ 0.265987f
C1205 a_3983_5056# _060_ 0.236911f
C1206 a_6003_10089# VPWR 0.221204f
C1207 _052_ _080_ 0.133809f
C1208 a_6982_4511# VPWR 0.199029f
C1209 ones[7] _049_ 0.108586f
C1210 clknet_1_0__leaf_clk a_1775_7125# 0.230932f
C1211 _091_ _011_ 0.28255f
C1212 _034_ counter\[9\] 0.965806f
C1213 _066_ net2 0.287208f
C1214 _077_ _047_ 1.19063f
C1215 net7 counter\[3\] 0.394746f
C1216 net9 a_1991_7691# 0.128527f
C1217 _050_ _049_ 0.406487f
C1218 _034_ _067_ 0.159912f
C1219 net1 clknet_1_1__leaf_clk 0.164762f
C1220 clknet_1_0__leaf_clk a_4227_2197# 0.236713f
C1221 _016_ _028_ 0.133649f
C1222 net4 a_9687_10927# 0.191132f
C1223 _037_ _040_ 0.194191f
C1224 a_9687_10927# VPWR 0.266989f
C1225 _068_ _072_ 0.325304f
C1226 counter\[4\] counter\[5\] 0.834767f
C1227 net1 _093_ 0.109442f
C1228 net3 net8 0.267648f
C1229 clknet_1_0__leaf_clk net2 0.812777f
C1230 net12 counter\[7\] 0.190311f
C1231 _050_ _052_ 0.3489f
C1232 _054_ clknet_0_clk 0.257127f
C1233 counter\[4\] _058_ 0.249037f
C1234 _063_ a_6633_5487# 0.253354f
C1235 net6 _071_ 0.1184f
C1236 net10 _024_ 0.246347f
C1237 net3 _034_ 0.180253f
C1238 a_8650_6153# _082_ 0.447234f
C1239 ones[1] _008_ 0.138855f
C1240 _070_ _080_ 0.14557f
C1241 a_1959_4949# a_2398_4943# 0.260055f
C1242 _086_ _057_ 0.113627f
C1243 net3 _088_ 0.246902f
C1244 net14 _022_ 0.899881f
C1245 a_3187_2251# _068_ 0.200381f
C1246 _000_ _084_ 0.224448f
C1247 _023_ a_4981_9991# 0.106529f
C1248 _036_ _035_ 0.451542f
C1249 a_3675_10601# a_3882_10660# 0.273138f
C1250 a_2807_7093# net10 0.128556f
C1251 net14 counter\[2\] 0.107472f
C1252 a_7171_10601# counter\[10\] 0.42622f
C1253 counter\[4\] _069_ 0.361285f
C1254 a_7001_8751# a_7442_8863# 0.110715f
C1255 _005_ a_7178_10505# 0.254948f
C1256 _090_ counter\[1\] 0.844393f
C1257 net6 _023_ 0.571739f
C1258 a_8999_6727# a_9095_6549# 0.310858f
C1259 net7 _001_ 1.09894f
C1260 a_3686_2767# a_3247_2773# 0.260055f
C1261 _023_ _036_ 0.144339f
C1262 counter\[1\] counter\[8\] 0.865566f
C1263 a_9933_5487# _004_ 0.131443f
C1264 _044_ _053_ 0.278679f
C1265 _049_ _047_ 0.184244f
C1266 _078_ _030_ 0.922502f
C1267 _068_ _052_ 0.177462f
C1268 _080_ net8 0.252063f
C1269 _005_ _068_ 0.116028f
C1270 _055_ VPWR 3.61182f
C1271 a_8643_6249# a_8650_6153# 0.959361f
C1272 net1 clknet_0_clk 0.277172f
C1273 _028_ _078_ 0.869744f
C1274 a_8650_6153# VPWR 0.272792f
C1275 net6 counter\[1\] 0.371854f
C1276 clknet_1_0__leaf_clk counter\[0\] 0.101026f
C1277 net1 _063_ 0.347892f
C1278 _038_ VPWR 1.56412f
C1279 _039_ counter\[1\] 0.558327f
C1280 _068_ _062_ 0.162107f
C1281 a_6173_3311# a_6871_3677# 0.191992f
C1282 net3 _028_ 0.104786f
C1283 a_6541_4399# counter\[3\] 0.32335f
C1284 _018_ _067_ 1.92125f
C1285 _048_ clknet_1_1__leaf_clk 0.136706f
C1286 net3 _091_ 0.442797f
C1287 ones[6] _054_ 0.14224f
C1288 a_6814_6031# VPWR 0.249185f
C1289 _088_ _080_ 0.425848f
C1290 _011_ VPWR 0.508466f
C1291 _009_ VPWR 0.609328f
C1292 a_8650_6153# a_8779_6409# 0.110715f
C1293 a_6982_4511# a_6814_4765# 0.239923f
C1294 a_9739_6005# VPWR 0.146462f
C1295 a_5399_3677# VPWR 0.179929f
C1296 _062_ _047_ 0.326709f
C1297 _079_ _026_ 0.100288f
C1298 _060_ _042_ 0.275542f
C1299 _025_ _087_ 0.144577f
C1300 net7 net12 0.332666f
C1301 a_6982_6005# a_6814_6031# 0.239923f
C1302 a_10239_9839# VPWR 0.263329f
C1303 _012_ VPWR 0.480176f
C1304 _063_ _033_ 0.200035f
C1305 counter\[2\] clknet_1_1__leaf_clk 0.208533f
C1306 _020_ _006_ 0.187493f
C1307 a_6887_10615# VPWR 0.226517f
C1308 _016_ VPWR 0.681845f
C1309 ones[3] net8 0.204655f
C1310 clknet_1_0__leaf_clk _084_ 0.187497f
C1311 _037_ _093_ 0.151362f
C1312 counter\[5\] net12 0.139738f
C1313 ones[7] a_7847_3855# 0.116737f
C1314 a_6007_3311# net4 0.109163f
C1315 _068_ _070_ 0.210377f
C1316 a_1941_7125# a_2639_7119# 0.194892f
C1317 a_6007_3311# VPWR 0.480261f
C1318 _038_ _015_ 0.319606f
C1319 a_8907_2986# _085_ 0.215739f
C1320 _081_ a_3797_6147# 0.205149f
C1321 clknet_1_0__leaf_clk a_4535_3311# 0.324838f
C1322 clknet_1_0__leaf_clk a_2111_6549# 0.28569f
C1323 net12 net9 0.134411f
C1324 pulse a_10199_3285# 0.237691f
C1325 _021_ _071_ 0.282492f
C1326 counter\[2\] a_7111_4221# 0.130274f
C1327 _058_ net12 0.271201f
C1328 _077_ net9 0.113841f
C1329 a_4974_3677# a_4535_3311# 0.260055f
C1330 net10 a_8459_4551# 0.171433f
C1331 a_9095_5461# VPWR 0.175438f
C1332 _068_ _031_ 0.14035f
C1333 a_7407_6005# counter\[1\] 0.130026f
C1334 _085_ net11 0.147729f
C1335 _078_ _082_ 0.16843f
C1336 _035_ _021_ 0.128593f
C1337 _062_ _087_ 0.220916f
C1338 counter\[9\] VPWR 2.87281f
C1339 _076_ a_9921_3476# 0.195965f
C1340 a_6719_10615# a_6887_10615# 0.310858f
C1341 a_8951_4949# _016_ 0.125574f
C1342 _086_ _024_ 0.372491f
C1343 counter\[4\] _079_ 0.184565f
C1344 _079_ a_9091_8439# 0.142329f
C1345 net14 _000_ 0.382458f
C1346 net7 a_7663_7485# 0.198783f
C1347 a_7274_9117# VPWR 0.258553f
C1348 a_6375_6037# a_6814_6031# 0.259379f
C1349 _013_ _037_ 0.356676f
C1350 _067_ VPWR 2.12863f
C1351 net5 _024_ 0.280592f
C1352 net12 a_7499_5755# 0.177551f
C1353 a_5843_4667# VPWR 0.432066f
C1354 _018_ _080_ 1.73097f
C1355 _005_ ones[0] 0.1221f
C1356 a_2971_8751# VPWR 0.481555f
C1357 net12 _056_ 0.168844f
C1358 a_6703_2197# VPWR 0.189881f
C1359 a_9558_4917# a_9117_4949# 0.110715f
C1360 _078_ VPWR 0.762695f
C1361 a_5960_5175# _068_ 0.15863f
C1362 a_8447_5175# _047_ 0.215864f
C1363 a_7407_4667# VPWR 0.437987f
C1364 counter\[6\] _078_ 0.120469f
C1365 _048_ a_6007_8207# 0.19449f
C1366 a_6169_6549# _053_ 0.137535f
C1367 counter\[5\] _049_ 0.208009f
C1368 _020_ _037_ 0.275821f
C1369 a_8999_5639# a_9095_5461# 0.310858f
C1370 net3 VPWR 5.02161f
C1371 a_2866_3087# _035_ 0.123674f
C1372 _043_ _042_ 0.250574f
C1373 net2 net11 0.785584f
C1374 a_2866_3087# _023_ 0.113501f
C1375 a_6423_11079# VPWR 0.200963f
C1376 _054_ _010_ 0.133437f
C1377 a_9213_3463# counter\[0\] 0.144163f
C1378 net1 a_8215_3861# 0.112696f
C1379 counter\[2\] counter\[10\] 0.2325f
C1380 _075_ VPWR 0.996037f
C1381 net1 counter\[1\] 0.285163f
C1382 counter\[10\] a_9435_9001# 0.109755f
C1383 _005_ net9 1.18715f
C1384 a_3973_7119# _043_ 0.11826f
C1385 _069_ _049_ 0.498793f
C1386 counter\[5\] _062_ 0.366672f
C1387 net2 _085_ 0.306726f
C1388 clknet_1_0__leaf_clk net14 0.627934f
C1389 _029_ _026_ 0.886961f
C1390 _028_ _047_ 0.123354f
C1391 _027_ _080_ 0.235157f
C1392 _091_ _047_ 0.231613f
C1393 _026_ _042_ 0.187765f
C1394 _080_ VPWR 6.62504f
C1395 clknet_1_0__leaf_clk net5 0.219217f
C1396 net6 _009_ 0.340088f
C1397 _019_ _029_ 1.04045f
C1398 a_7442_8863# a_7274_9117# 0.239923f
C1399 a_6729_6031# _001_ 0.114649f
C1400 _006_ counter\[1\] 0.621884f
C1401 a_8907_2986# _008_ 0.130228f
C1402 _018_ _068_ 2.42344f
C1403 ones[0] net8 0.141717f
C1404 _023_ _081_ 0.251007f
C1405 a_3811_10761# a_3675_10601# 0.141453f
C1406 _033_ counter\[1\] 0.102013f
C1407 counter\[0\] net11 0.181537f
C1408 a_9091_10004# _067_ 0.189198f
C1409 a_10287_6250# _082_ 0.219149f
C1410 a_7378_10660# VPWR 0.25986f
C1411 counter\[3\] _060_ 0.157965f
C1412 ones[2] net13 0.197794f
C1413 _077_ _079_ 0.128829f
C1414 _039_ _012_ 0.180951f
C1415 net7 _031_ 0.112093f
C1416 a_4627_5056# VPWR 0.186843f
C1417 counter\[4\] _060_ 0.350954f
C1418 _060_ a_9091_8439# 0.171617f
C1419 _076_ counter\[4\] 0.123928f
C1420 ones[7] VPWR 0.410013f
C1421 a_9079_3855# a_8381_3861# 0.191992f
C1422 a_2125_4949# a_2823_4943# 0.192206f
C1423 counter\[7\] _091_ 1.72702f
C1424 a_6835_8751# VPWR 0.48298f
C1425 _088_ a_3847_8903# 0.201282f
C1426 _022_ _071_ 0.161448f
C1427 a_10239_7663# VPWR 0.21428f
C1428 _066_ _059_ 0.163455f
C1429 a_4731_4233# VPWR 0.173905f
C1430 a_6927_9301# a_7093_9301# 0.961627f
C1431 _037_ _071_ 0.579837f
C1432 counter\[4\] _029_ 0.259824f
C1433 net7 net8 0.224932f
C1434 _037_ a_6283_7669# 0.156226f
C1435 a_9871_2223# VPWR 0.231477f
C1436 counter\[9\] counter\[8\] 0.195261f
C1437 a_8390_7119# VPWR 1.372f
C1438 a_9379_5461# _004_ 0.117471f
C1439 _050_ VPWR 1.9988f
C1440 counter\[3\] _042_ 1.12298f
C1441 a_10147_4399# net14 0.188603f
C1442 _010_ _006_ 0.141203f
C1443 a_3431_4943# _060_ 0.100183f
C1444 net9 _031_ 0.494815f
C1445 net10 net11 1.16302f
C1446 ones[3] VPWR 0.455781f
C1447 _085_ _008_ 0.140535f
C1448 counter\[5\] net8 0.111447f
C1449 a_10287_6250# VPWR 0.256423f
C1450 _020_ _024_ 0.534392f
C1451 a_7123_2223# a_6987_2197# 0.136009f
C1452 a_4535_3311# _074_ 0.435294f
C1453 net6 counter\[9\] 0.105953f
C1454 a_9919_4087# _026_ 0.226924f
C1455 net9 net8 1.59469f
C1456 a_1499_5056# VPWR 0.238377f
C1457 clknet_1_0__leaf_clk _059_ 0.312591f
C1458 a_7178_10505# VPWR 0.327826f
C1459 a_5507_10357# net3 0.123754f
C1460 _043_ _026_ 0.133137f
C1461 a_6173_3311# _074_ 0.466737f
C1462 a_9739_6005# a_9915_6337# 0.185422f
C1463 a_5960_5175# a_5687_5175# 0.167615f
C1464 _090_ net3 0.177894f
C1465 net6 a_2971_8751# 0.254897f
C1466 a_7074_5599# VPWR 0.193161f
C1467 net3 counter\[8\] 0.109785f
C1468 _068_ VPWR 3.25522f
C1469 counter\[2\] counter\[1\] 2.07228f
C1470 _078_ _039_ 0.191528f
C1471 net6 net3 0.488668f
C1472 _047_ VPWR 3.56807f
C1473 _021_ _009_ 0.747461f
C1474 net3 _036_ 0.156612f
C1475 _043_ a_1941_7125# 0.458765f
C1476 _054_ a_9739_6005# 0.113498f
C1477 _074_ a_4668_7913# 0.100587f
C1478 net7 _014_ 0.829201f
C1479 net2 _008_ 0.414302f
C1480 net7 _028_ 0.523386f
C1481 _053_ clknet_0_clk 0.382571f
C1482 clknet_1_0__leaf_clk clknet_0_clk 0.216514f
C1483 a_7442_8863# a_6835_8751# 0.136009f
C1484 a_7001_8751# _022_ 0.180977f
C1485 ready a_10147_4399# 0.109593f
C1486 counter\[2\] _010_ 0.138341f
C1487 counter\[5\] _091_ 0.129362f
C1488 net6 _075_ 0.131895f
C1489 _019_ _026_ 0.167568f
C1490 _010_ a_9435_9001# 0.106246f
C1491 a_6475_7913# _031_ 0.154609f
C1492 a_6987_2197# VPWR 0.404043f
C1493 _068_ _015_ 0.685636f
C1494 _066_ counter\[10\] 0.115793f
C1495 a_7980_4649# _030_ 0.10606f
C1496 counter\[7\] net4 0.211439f
C1497 _020_ _053_ 0.181925f
C1498 a_3247_2773# VPWR 0.438154f
C1499 _056_ a_2191_10615# 0.141633f
C1500 clknet_1_0__leaf_clk _020_ 0.331268f
C1501 counter\[7\] VPWR 1.23693f
C1502 _028_ net9 0.584181f
C1503 _055_ net13 0.501995f
C1504 _077_ _060_ 0.448252f
C1505 _080_ counter\[8\] 0.281898f
C1506 a_4811_4399# VPWR 0.685681f
C1507 _045_ _040_ 0.338469f
C1508 _028_ _041_ 0.119878f
C1509 net2 net10 0.39543f
C1510 _058_ _091_ 0.132367f
C1511 a_7331_5853# a_7499_5755# 0.310858f
C1512 a_3983_5056# _062_ 0.124043f
C1513 a_4535_7232# VPWR 0.201534f
C1514 net2 _084_ 0.135956f
C1515 counter\[6\] counter\[7\] 0.620944f
C1516 a_7847_3133# VPWR 0.408571f
C1517 net1 _011_ 0.600464f
C1518 _087_ VPWR 4.06231f
C1519 net14 _083_ 0.214398f
C1520 net6 _080_ 0.647339f
C1521 counter\[5\] _018_ 0.431767f
C1522 a_4311_4087# VPWR 0.191489f
C1523 net12 _042_ 0.425247f
C1524 counter\[3\] _026_ 0.236759f
C1525 a_2214_7119# VPWR 0.274883f
C1526 _052_ _003_ 0.100156f
C1527 _069_ _091_ 0.631932f
C1528 _086_ _074_ 0.206343f
C1529 _023_ _024_ 0.73084f
C1530 net14 net11 0.118267f
C1531 _033_ _038_ 0.220806f
C1532 net1 _016_ 0.337872f
C1533 a_7699_9117# VPWR 0.196304f
C1534 _044_ net10 0.405106f
C1535 a_3847_8903# VPWR 0.215427f
C1536 _013_ a_4781_2223# 0.114651f
C1537 a_8999_6727# VPWR 0.393393f
C1538 _045_ net5 0.226994f
C1539 ones[0] VPWR 0.293252f
C1540 net6 a_9871_2223# 0.19921f
C1541 net6 _050_ 3.05294f
C1542 net14 _085_ 0.410451f
C1543 _039_ a_8390_7119# 0.110278f
C1544 a_3697_6031# VPWR 0.167969f
C1545 _092_ _060_ 0.195801f
C1546 _004_ clknet_1_1__leaf_clk 0.858585f
C1547 a_6519_9813# a_6810_10113# 0.192341f
C1548 a_7867_9019# a_7699_9117# 0.310858f
C1549 _058_ _082_ 1.73234f
C1550 _084_ _008_ 0.21741f
C1551 net1 counter\[9\] 0.127843f
C1552 _005_ a_3682_10505# 0.258403f
C1553 a_3811_10761# a_3882_10660# 0.239923f
C1554 counter\[1\] _073_ 0.160215f
C1555 a_6803_9813# a_6939_9839# 0.136009f
C1556 a_6810_10113# _008_ 0.180977f
C1557 a_4227_2197# a_4363_2223# 0.141453f
C1558 a_5843_4667# a_5675_4765# 0.310858f
C1559 net7 net4 0.107977f
C1560 _003_ _070_ 5.74987f
C1561 _002_ VPWR 1.357f
C1562 net7 VPWR 5.20652f
C1563 _068_ counter\[8\] 2.9687f
C1564 _000_ a_4627_6031# 0.109291f
C1565 a_5687_5175# VPWR 0.194149f
C1566 net2 _040_ 0.312982f
C1567 a_6982_4511# a_6375_4399# 0.136009f
C1568 net1 a_2971_8751# 0.129992f
C1569 _043_ net12 0.688549f
C1570 net7 counter\[6\] 0.104914f
C1571 a_5142_3423# VPWR 0.177211f
C1572 counter\[5\] VPWR 1.63816f
C1573 a_6703_2197# a_6994_2497# 0.194215f
C1574 _061_ a_4627_6031# 0.193133f
C1575 _067_ net13 0.889293f
C1576 net1 _078_ 0.885598f
C1577 net6 _068_ 0.956181f
C1578 a_6515_4074# VPWR 0.255101f
C1579 clknet_1_0__leaf_clk _035_ 0.109685f
C1580 counter\[6\] counter\[5\] 0.337916f
C1581 net9 VPWR 3.79191f
C1582 _062_ _060_ 0.358295f
C1583 _076_ _062_ 0.183961f
C1584 a_7980_4649# VPWR 0.153671f
C1585 _058_ VPWR 1.53159f
C1586 _059_ net11 0.741368f
C1587 _041_ VPWR 0.463551f
C1588 a_4802_4132# a_4731_4233# 0.239923f
C1589 a_2111_6549# net10 0.148574f
C1590 clknet_1_0__leaf_clk _023_ 1.39567f
C1591 a_7407_4667# a_7239_4765# 0.310858f
C1592 net1 net3 0.782649f
C1593 a_3686_2767# a_3854_2741# 0.239923f
C1594 net6 _047_ 0.106143f
C1595 a_5399_3677# a_4701_3311# 0.190502f
C1596 a_7886_3311# _028_ 0.113303f
C1597 a_7171_10601# a_7378_10660# 0.260055f
C1598 net14 net2 0.604967f
C1599 net3 net13 0.132691f
C1600 a_9213_3463# _063_ 0.10606f
C1601 _064_ _060_ 0.100706f
C1602 a_2665_6575# _009_ 0.114646f
C1603 _069_ VPWR 2.56134f
C1604 a_3391_10615# VPWR 0.197955f
C1605 _090_ _087_ 0.125216f
C1606 a_7499_5755# VPWR 0.431814f
C1607 _076_ _070_ 0.182592f
C1608 a_8631_2986# _014_ 0.110677f
C1609 a_6927_9301# a_7366_9295# 0.260055f
C1610 _056_ VPWR 1.69189f
C1611 a_2409_4445# VPWR 0.160428f
C1612 a_9379_6549# a_9586_6549# 0.273138f
C1613 a_9386_6849# a_9515_6575# 0.111047f
C1614 _043_ _025_ 0.526977f
C1615 _020_ _083_ 0.352066f
C1616 clknet_0_clk net11 0.167732f
C1617 _005_ a_9921_3476# 0.130271f
C1618 _057_ counter\[9\] 0.140858f
C1619 net3 _081_ 0.112013f
C1620 a_7171_10601# a_7178_10505# 0.96403f
C1621 _063_ net11 0.184628f
C1622 _039_ _087_ 0.194442f
C1623 _029_ _031_ 0.127825f
C1624 a_9091_10004# _002_ 0.108492f
C1625 _060_ net8 0.317157f
C1626 a_7281_9295# _012_ 0.128307f
C1627 _080_ net13 0.194409f
C1628 a_2697_2767# VPWR 0.220144f
C1629 a_6541_4399# VPWR 0.300619f
C1630 net14 counter\[0\] 0.658249f
C1631 counter\[2\] counter\[9\] 0.459245f
C1632 _014_ _003_ 0.195926f
C1633 _040_ net10 0.121543f
C1634 clk _025_ 0.250006f
C1635 _086_ counter\[0\] 1.25671f
C1636 pulse _005_ 0.128656f
C1637 counter\[4\] net12 0.186252f
C1638 a_6475_7913# VPWR 0.119909f
C1639 a_4345_6031# _092_ 0.144594f
C1640 counter\[4\] _077_ 0.178138f
C1641 _034_ _060_ 0.321664f
C1642 _081_ _075_ 0.138526f
C1643 a_1460_9269# VPWR 0.266812f
C1644 net5 counter\[0\] 0.585088f
C1645 a_6425_10602# _018_ 0.131141f
C1646 _093_ net2 0.218195f
C1647 a_6633_5487# a_7074_5599# 0.110715f
C1648 _088_ _060_ 0.605591f
C1649 a_10239_10383# net8 0.211204f
C1650 a_5418_4511# VPWR 0.179436f
C1651 _025_ _026_ 0.404821f
C1652 net7 a_5507_10357# 0.173021f
C1653 a_4521_8903# net2 0.111974f
C1654 clk _052_ 0.2701f
C1655 _045_ counter\[10\] 0.309915f
C1656 _018_ _003_ 0.115507f
C1657 _034_ _042_ 0.361691f
C1658 a_4602_3977# VPWR 0.28554f
C1659 a_9558_4917# VPWR 0.183851f
C1660 _050_ net13 0.17173f
C1661 net14 _084_ 0.240691f
C1662 _086_ net10 0.102977f
C1663 a_2639_7119# VPWR 0.197803f
C1664 net3 counter\[2\] 0.734566f
C1665 a_4697_5461# VPWR 1.19839f
C1666 _086_ _084_ 0.110315f
C1667 counter\[4\] _072_ 0.139215f
C1668 rst a_10199_2197# 0.244783f
C1669 _013_ a_4227_2197# 0.100274f
C1670 a_7886_3311# VPWR 0.459947f
C1671 _044_ clknet_1_1__leaf_clk 0.370847f
C1672 net5 net10 0.147308f
C1673 a_5141_4917# _075_ 0.114629f
C1674 _050_ _006_ 0.897976f
C1675 a_2460_3971# _088_ 0.111265f
C1676 _079_ VPWR 0.297085f
C1677 net7 _039_ 0.409923f
C1678 _012_ _024_ 0.1749f
C1679 a_10147_4399# _051_ 0.122182f
C1680 _014_ _060_ 0.230092f
C1681 counter\[0\] clknet_1_1__leaf_clk 0.578338f
C1682 _076_ _028_ 0.753369f
C1683 a_6541_6037# a_7239_6031# 0.194215f
C1684 net14 _032_ 0.120635f
C1685 _008_ clknet_1_1__leaf_clk 0.376466f
C1686 a_3983_5056# VPWR 0.204957f
C1687 _054_ counter\[7\] 0.184644f
C1688 a_8631_2986# VPWR 0.194085f
C1689 a_4234_2497# a_3943_2197# 0.194892f
C1690 net2 a_10199_2197# 0.17126f
C1691 counter\[4\] _025_ 0.143749f
C1692 a_9558_4917# a_8951_4949# 0.141453f
C1693 _057_ _080_ 0.13119f
C1694 counter\[0\] a_7111_4221# 0.150439f
C1695 a_9919_4087# net8 0.27724f
C1696 _042_ _030_ 0.235237f
C1697 ready _008_ 0.169188f
C1698 _074_ _071_ 0.424511f
C1699 a_2555_10704# a_2191_10615# 0.124682f
C1700 _073_ _012_ 0.440412f
C1701 _041_ _039_ 0.271276f
C1702 a_2682_3311# VPWR 0.200511f
C1703 a_1731_6727# VPWR 0.435673f
C1704 _028_ _042_ 0.105118f
C1705 _020_ net2 0.102998f
C1706 a_7378_10660# a_7307_10761# 0.239923f
C1707 a_6425_10602# VPWR 0.231425f
C1708 a_5717_4087# _080_ 0.116814f
C1709 a_9213_3463# counter\[1\] 0.216311f
C1710 net10 clknet_1_1__leaf_clk 0.194854f
C1711 counter\[9\] _024_ 0.632698f
C1712 _033_ _068_ 0.112334f
C1713 _023_ _074_ 0.231249f
C1714 _003_ net4 0.225347f
C1715 a_8256_11177# _068_ 0.104274f
C1716 _003_ VPWR 2.84873f
C1717 a_6810_10113# clknet_1_1__leaf_clk 0.311852f
C1718 _038_ _053_ 0.110413f
C1719 a_5567_3579# VPWR 0.403151f
C1720 a_6994_2497# a_6987_2197# 0.962054f
C1721 _059_ net10 0.132151f
C1722 _044_ clknet_0_clk 0.484879f
C1723 _026_ _031_ 0.578228f
C1724 _023_ _045_ 0.112385f
C1725 a_9379_5461# clknet_1_1__leaf_clk 0.320537f
C1726 clknet_1_0__leaf_clk _011_ 0.690835f
C1727 counter\[9\] _073_ 0.376501f
C1728 a_9096_4373# VPWR 0.16185f
C1729 a_10199_3285# VPWR 0.357209f
C1730 clknet_1_0__leaf_clk _009_ 0.183204f
C1731 _026_ net8 0.277476f
C1732 net1 _087_ 0.402916f
C1733 counter\[1\] net11 0.524259f
C1734 a_7178_10505# a_7307_10761# 0.118966f
C1735 _010_ _004_ 0.84686f
C1736 net3 _024_ 0.353322f
C1737 a_6927_9301# VPWR 0.479911f
C1738 counter\[9\] _017_ 0.591276f
C1739 a_8109_5639# net11 0.171766f
C1740 _019_ net8 0.231126f
C1741 _059_ _089_ 0.33475f
C1742 _078_ _073_ 0.321067f
C1743 clknet_1_0__leaf_clk a_6007_3311# 0.214796f
C1744 _043_ _030_ 0.218824f
C1745 counter\[4\] _070_ 0.352217f
C1746 _066_ counter\[9\] 0.440752f
C1747 a_6541_6037# clknet_1_1__leaf_clk 0.112405f
C1748 a_3682_10505# VPWR 0.302578f
C1749 _088_ _026_ 0.220282f
C1750 a_9586_6549# VPWR 0.251851f
C1751 net7 _054_ 0.227138f
C1752 _006_ _087_ 0.61736f
C1753 a_4215_4087# a_4311_4087# 0.310858f
C1754 a_9379_5461# a_9515_5487# 0.141453f
C1755 net3 _061_ 0.325793f
C1756 _057_ _068_ 0.185231f
C1757 a_1991_7691# net8 0.16196f
C1758 a_4234_2497# VPWR 0.29986f
C1759 net3 _073_ 0.134907f
C1760 _048_ _047_ 0.222836f
C1761 counter\[7\] _081_ 0.102214f
C1762 _060_ VPWR 5.77302f
C1763 a_2382_7093# a_2214_7119# 0.239923f
C1764 _076_ VPWR 0.849015f
C1765 _037_ _068_ 0.352388f
C1766 _063_ _084_ 0.296982f
C1767 counter\[2\] _068_ 0.152309f
C1768 _000_ _075_ 0.246839f
C1769 _029_ _027_ 0.820087f
C1770 _076_ counter\[6\] 0.248311f
C1771 clknet_1_0__leaf_clk counter\[9\] 0.92438f
C1772 _058_ _054_ 0.144399f
C1773 a_4580_8439# VPWR 0.170199f
C1774 _029_ VPWR 0.948896f
C1775 _090_ _079_ 0.30763f
C1776 a_6607_2375# VPWR 0.390429f
C1777 _042_ VPWR 1.4468f
C1778 _066_ net3 0.335488f
C1779 a_10239_10383# VPWR 0.250065f
C1780 _032_ clknet_0_clk 0.206539f
C1781 _014_ _026_ 0.314891f
C1782 _005_ a_4229_10761# 0.114823f
C1783 net1 net7 1.21551f
C1784 _028_ _026_ 0.252715f
C1785 counter\[3\] a_2191_10615# 0.166583f
C1786 net12 _052_ 0.114042f
C1787 counter\[6\] _042_ 0.739724f
C1788 ones[10] VPWR 0.352948f
C1789 counter\[10\] _084_ 0.124988f
C1790 a_2460_3971# VPWR 0.16886f
C1791 net7 net13 0.480774f
C1792 a_7074_5599# a_6906_5853# 0.239923f
C1793 a_9832_8181# _069_ 0.111658f
C1794 _076_ _015_ 0.176272f
C1795 net14 clknet_1_1__leaf_clk 0.188082f
C1796 a_3973_7119# VPWR 0.181274f
C1797 a_5149_4233# _020_ 0.125406f
C1798 clknet_1_0__leaf_clk net3 0.110525f
C1799 rst ones[2] 0.242446f
C1800 a_7039_3579# counter\[3\] 0.126181f
C1801 _037_ a_4535_7232# 0.216004f
C1802 _043_ _082_ 0.200578f
C1803 a_6423_9991# VPWR 0.407894f
C1804 a_9983_4917# VPWR 0.406328f
C1805 net5 clknet_1_1__leaf_clk 0.781304f
C1806 a_2555_10704# VPWR 0.239642f
C1807 net14 a_4521_8903# 0.17326f
C1808 a_4580_8439# a_4307_8439# 0.167615f
C1809 net5 _093_ 0.710202f
C1810 a_6939_9839# VPWR 0.196209f
C1811 a_6169_6549# clknet_0_clk 1.72801f
C1812 a_4595_4073# a_4731_4233# 0.136009f
C1813 _086_ a_1683_10496# 0.154223f
C1814 a_9435_9001# _087_ 0.111073f
C1815 a_9921_3476# VPWR 0.20838f
C1816 _028_ counter\[3\] 0.14579f
C1817 _066_ _080_ 0.124025f
C1818 net5 _059_ 0.615846f
C1819 clknet_1_0__leaf_clk _075_ 0.116451f
C1820 net9 _006_ 0.443036f
C1821 counter\[4\] _028_ 0.95183f
C1822 ones[5] VPWR 0.323968f
C1823 ones[2] net2 0.328529f
C1824 a_3854_2741# VPWR 0.196357f
C1825 a_8175_6549# _025_ 0.17201f
C1826 _033_ net9 0.335078f
C1827 a_9919_4087# VPWR 0.206425f
C1828 a_2318_6549# VPWR 0.268796f
C1829 a_10239_7663# ones[1] 0.114396f
C1830 _043_ _027_ 0.356343f
C1831 _043_ net4 0.342651f
C1832 _044_ counter\[1\] 0.10346f
C1833 pulse VPWR 0.119216f
C1834 _043_ VPWR 1.60634f
C1835 _055_ _074_ 0.270272f
C1836 a_2318_6549# a_2247_6575# 0.239923f
C1837 a_9386_6849# clknet_1_1__leaf_clk 0.369315f
C1838 ones[3] ones[1] 0.103553f
C1839 clknet_1_0__leaf_clk _080_ 1.30193f
C1840 _018_ counter\[3\] 0.489367f
C1841 _044_ a_8109_5639# 0.106013f
C1842 counter\[0\] counter\[1\] 3.83085f
C1843 a_2513_3561# VPWR 0.266861f
C1844 a_2118_6849# VPWR 0.352571f
C1845 net7 _048_ 0.148342f
C1846 _065_ VPWR 1.75159f
C1847 clk VPWR 0.633935f
C1848 net12 net8 0.10463f
C1849 _038_ net11 0.141591f
C1850 _077_ net8 0.101169f
C1851 _062_ _049_ 0.110331f
C1852 a_4345_6031# VPWR 0.162465f
C1853 a_9386_5761# VPWR 0.303643f
C1854 _065_ counter\[6\] 0.609724f
C1855 a_2247_6575# a_2118_6849# 0.110715f
C1856 net14 _020_ 0.623777f
C1857 _034_ net12 0.278941f
C1858 _026_ _027_ 1.19555f
C1859 a_7239_4765# a_6541_4399# 0.192016f
C1860 net7 _037_ 0.442569f
C1861 _060_ counter\[8\] 0.237623f
C1862 a_5141_4917# counter\[5\] 0.217876f
C1863 a_4123_9514# VPWR 0.275888f
C1864 _026_ VPWR 2.69971f
C1865 a_6987_2197# a_7194_2197# 0.260055f
C1866 net7 counter\[2\] 0.113593f
C1867 a_4701_3311# a_5142_3423# 0.110672f
C1868 a_3799_10927# _060_ 0.165768f
C1869 net5 _020_ 0.115804f
C1870 _005_ _062_ 0.20806f
C1871 counter\[1\] net10 0.145079f
C1872 a_2509_4663# _075_ 0.203874f
C1873 a_8381_3861# a_8215_3861# 0.970499f
C1874 _084_ counter\[1\] 0.377432f
C1875 net6 _060_ 1.04693f
C1876 a_5165_4399# _000_ 0.113524f
C1877 net14 counter\[10\] 0.219716f
C1878 _019_ VPWR 0.734878f
C1879 a_6007_3311# _074_ 0.100377f
C1880 a_4811_4399# a_4977_4399# 0.966391f
C1881 _037_ net9 0.136882f
C1882 _039_ _060_ 1.74184f
C1883 a_1679_10089# VPWR 0.237684f
C1884 counter\[2\] net9 0.291939f
C1885 a_7357_9839# _008_ 0.114644f
C1886 _037_ _041_ 0.333063f
C1887 _019_ a_6821_5487# 0.120224f
C1888 _046_ _032_ 0.585833f
C1889 a_1991_7691# VPWR 0.244385f
C1890 ones[10] counter\[8\] 0.13881f
C1891 _051_ _008_ 1.09577f
C1892 a_3029_6031# VPWR 0.193358f
C1893 a_1941_7125# VPWR 0.358133f
C1894 _083_ counter\[9\] 0.173161f
C1895 a_5087_6575# VPWR 0.217457f
C1896 clknet_0_clk clknet_1_1__leaf_clk 0.121177f
C1897 counter\[3\] net4 0.688758f
C1898 ones[2] _084_ 0.372937f
C1899 _052_ _070_ 1.96964f
C1900 _039_ _042_ 0.117139f
C1901 net12 _030_ 0.466567f
C1902 _007_ VPWR 0.38574f
C1903 counter\[3\] VPWR 2.71991f
C1904 a_2566_4917# VPWR 0.195559f
C1905 _074_ counter\[9\] 0.579438f
C1906 _063_ clknet_1_1__leaf_clk 0.256375f
C1907 counter\[4\] net4 0.478066f
C1908 _010_ _084_ 0.25354f
C1909 _069_ counter\[2\] 0.3375f
C1910 _028_ net12 0.364498f
C1911 clknet_1_0__leaf_clk _068_ 0.118245f
C1912 _057_ _056_ 0.168777f
C1913 a_4434_2197# VPWR 0.253146f
C1914 counter\[4\] VPWR 3.15271f
C1915 a_9091_8439# VPWR 0.203595f
C1916 _028_ _077_ 0.381764f
C1917 _020_ clknet_1_1__leaf_clk 0.174193f
C1918 _005_ _031_ 0.913695f
C1919 _020_ _093_ 0.147905f
C1920 _053_ _047_ 0.283983f
C1921 a_7886_3311# _033_ 0.160941f
C1922 a_3431_4943# VPWR 0.194787f
C1923 _052_ net8 0.114831f
C1924 _005_ net8 1.21343f
C1925 counter\[10\] clknet_1_1__leaf_clk 0.397211f
C1926 _074_ net3 0.110877f
C1927 counter\[3\] _015_ 0.21164f
C1928 _005_ _034_ 0.10791f
C1929 a_7093_9301# VPWR 0.291326f
C1930 a_9117_4949# VPWR 0.299238f
C1931 a_10195_7338# VPWR 0.23678f
C1932 clknet_1_0__leaf_clk a_3247_2773# 0.295647f
C1933 clknet_1_0__leaf_clk counter\[7\] 0.550674f
C1934 _045_ net3 0.447967f
C1935 _010_ a_10239_8751# 0.109783f
C1936 clknet_1_0__leaf_clk a_4811_4399# 0.292864f
C1937 _001_ VPWR 1.19845f
C1938 _003_ net13 0.106676f
C1939 net5 _035_ 0.453203f
C1940 counter\[4\] a_8999_5639# 0.129228f
C1941 _021_ _060_ 0.325845f
C1942 _076_ _021_ 0.245263f
C1943 a_7791_9295# a_7093_9301# 0.190773f
C1944 net1 a_9096_4373# 0.137342f
C1945 net1 a_10199_3285# 0.171313f
C1946 net5 a_7959_9269# 0.155412f
C1947 _023_ net5 1.17615f
C1948 _028_ _092_ 0.309502f
C1949 _028_ _049_ 0.129855f
C1950 _091_ _092_ 0.229005f
C1951 net14 counter\[1\] 0.630316f
C1952 counter\[0\] _038_ 0.416541f
C1953 _034_ _064_ 0.711015f
C1954 _044_ _009_ 0.332075f
C1955 net6 clk 0.109816f
C1956 a_2682_3311# _081_ 0.114442f
C1957 _086_ a_7419_5281# 0.158071f
C1958 a_9095_6549# VPWR 0.187925f
C1959 a_8951_4949# a_9117_4949# 0.969958f
C1960 counter\[0\] _011_ 0.232775f
C1961 net5 counter\[1\] 0.484273f
C1962 _080_ net11 1.19811f
C1963 _019_ counter\[8\] 0.155715f
C1964 _085_ _075_ 0.313092f
C1965 net12 net4 0.582357f
C1966 _036_ _026_ 0.1146f
C1967 _093_ _071_ 0.142749f
C1968 _039_ _026_ 0.191513f
C1969 net12 VPWR 4.41379f
C1970 _077_ VPWR 0.909885f
C1971 net1 _076_ 0.147769f
C1972 a_8822_3829# VPWR 0.181893f
C1973 _066_ counter\[5\] 0.291495f
C1974 net14 a_7001_8751# 0.45912f
C1975 _056_ _024_ 0.814662f
C1976 a_6803_9813# VPWR 0.462201f
C1977 a_6375_4399# a_6541_4399# 0.960208f
C1978 _060_ net13 0.395344f
C1979 _076_ net13 0.214701f
C1980 _034_ net8 0.332681f
C1981 _090_ counter\[3\] 1.39266f
C1982 _017_ _041_ 0.165828f
C1983 a_6375_6037# _001_ 0.120049f
C1984 a_5363_2880# _060_ 0.194155f
C1985 counter\[3\] counter\[8\] 0.118791f
C1986 _011_ _084_ 0.394972f
C1987 _009_ net10 0.124503f
C1988 a_6467_5487# a_7074_5599# 0.136009f
C1989 net6 a_3029_6031# 0.143138f
C1990 a_9586_5461# VPWR 0.250706f
C1991 _023_ _059_ 1.00803f
C1992 _028_ _064_ 0.131965f
C1993 clknet_1_0__leaf_clk net7 0.125697f
C1994 net3 net2 0.263692f
C1995 _050_ net11 0.196401f
C1996 a_8215_3861# clknet_1_1__leaf_clk 0.250105f
C1997 a_6614_3423# VPWR 0.178619f
C1998 _082_ _092_ 0.12393f
C1999 counter\[1\] clknet_1_1__leaf_clk 0.537122f
C2000 a_3686_2767# VPWR 0.259694f
C2001 clknet_1_0__leaf_clk counter\[5\] 0.690222f
C2002 _072_ VPWR 0.625834f
C2003 _076_ _033_ 0.206759f
C2004 _034_ _088_ 0.147721f
C2005 a_5142_3423# a_4974_3677# 0.239923f
C2006 a_1499_5056# _074_ 0.104745f
C2007 _033_ a_4580_8439# 0.120859f
C2008 a_8654_3855# a_8215_3861# 0.271965f
C2009 _043_ _021_ 0.358032f
C2010 a_7111_4221# counter\[1\] 0.15777f
C2011 clknet_1_0__leaf_clk _058_ 0.340444f
C2012 counter\[4\] _039_ 0.793323f
C2013 a_7663_7485# VPWR 0.415036f
C2014 ones[6] counter\[10\] 0.227739f
C2015 _054_ _043_ 0.862407f
C2016 _017_ _056_ 0.621392f
C2017 a_4977_4399# a_5418_4511# 0.110715f
C2018 a_4811_4399# a_5250_4765# 0.273138f
C2019 _067_ counter\[0\] 0.123175f
C2020 _081_ _060_ 0.356758f
C2021 _076_ _081_ 0.236153f
C2022 a_5843_4667# counter\[0\] 0.127039f
C2023 _033_ _042_ 0.133796f
C2024 a_3973_7119# a_4073_7235# 0.167615f
C2025 _025_ net4 0.126176f
C2026 _074_ _068_ 0.260831f
C2027 _025_ VPWR 0.618222f
C2028 _050_ a_9687_4399# 0.19771f
C2029 a_3187_2251# VPWR 0.225231f
C2030 counter\[0\] _078_ 0.167534f
C2031 _092_ VPWR 0.385388f
C2032 _018_ _070_ 0.20096f
C2033 _049_ VPWR 1.72413f
C2034 a_1867_4399# VPWR 0.252429f
C2035 a_8175_6549# VPWR 0.169677f
C2036 a_6173_3311# a_6007_3311# 0.963466f
C2037 net2 _080_ 0.669142f
C2038 net3 counter\[0\] 1.3442f
C2039 a_2991_4917# VPWR 0.421477f
C2040 a_8447_5175# _028_ 0.193558f
C2041 _018_ _031_ 0.115506f
C2042 _034_ _028_ 0.6722f
C2043 a_4595_4073# a_4602_3977# 0.959647f
C2044 _052_ net4 0.118859f
C2045 net3 _008_ 0.660796f
C2046 _021_ _026_ 0.276438f
C2047 _052_ VPWR 2.84138f
C2048 a_3413_2773# a_3247_2773# 0.959361f
C2049 _051_ _093_ 1.30587f
C2050 _005_ VPWR 1.76856f
C2051 a_8359_6263# a_8263_6263# 0.310858f
C2052 _054_ _026_ 0.138085f
C2053 a_7939_6031# VPWR 0.231635f
C2054 net1 _043_ 0.190058f
C2055 a_2807_7093# a_2639_7119# 0.310858f
C2056 _063_ counter\[1\] 0.664225f
C2057 _009_ _040_ 0.222622f
C2058 _019_ a_6633_5487# 0.247017f
C2059 _043_ net13 0.142394f
C2060 _062_ VPWR 1.08126f
C2061 a_9435_9001# _060_ 0.113164f
C2062 net1 clk 0.108291f
C2063 net3 net10 0.342531f
C2064 _086_ _055_ 2.20005f
C2065 _050_ net2 0.82616f
C2066 net3 _084_ 0.906939f
C2067 _079_ _073_ 0.107249f
C2068 clk net13 0.120993f
C2069 _037_ _042_ 0.289592f
C2070 _064_ VPWR 0.643632f
C2071 a_8447_8916# _079_ 0.180207f
C2072 _043_ _033_ 0.200322f
C2073 _028_ _030_ 0.533066f
C2074 _054_ a_5087_6575# 0.219023f
C2075 counter\[10\] counter\[1\] 0.108207f
C2076 _014_ _028_ 0.445124f
C2077 net5 _038_ 0.170342f
C2078 net1 _026_ 0.277587f
C2079 _028_ _091_ 0.470778f
C2080 _070_ VPWR 1.59632f
C2081 counter\[7\] _085_ 0.862816f
C2082 a_9832_8181# counter\[3\] 0.1869f
C2083 net12 _039_ 0.198966f
C2084 counter\[6\] _070_ 0.142035f
C2085 _034_ _082_ 0.103523f
C2086 net5 _009_ 0.12024f
C2087 clknet_1_0__leaf_clk a_4602_3977# 0.205456f
C2088 net3 _089_ 0.380056f
C2089 _017_ a_2129_7119# 0.131384f
C2090 _031_ VPWR 1.62615f
C2091 counter\[9\] _040_ 0.92302f
C2092 _068_ net2 0.281465f
C2093 a_2409_4445# a_2509_4663# 0.167615f
C2094 clknet_1_0__leaf_clk a_4697_5461# 1.80219f
C2095 net5 _012_ 0.419547f
C2096 _072_ counter\[8\] 1.65239f
C2097 _084_ _080_ 0.134257f
C2098 _033_ _026_ 0.567332f
C2099 a_9379_6549# VPWR 0.67138f
C2100 a_8447_8439# _028_ 0.201408f
C2101 _067_ _040_ 1.28885f
C2102 a_3799_10927# _072_ 0.209864f
C2103 net8 VPWR 2.45944f
C2104 a_7366_9295# VPWR 0.239492f
C2105 _043_ _048_ 0.234468f
C2106 _038_ clknet_1_1__leaf_clk 0.225012f
C2107 a_8447_5175# VPWR 0.200482f
C2108 _034_ VPWR 1.99971f
C2109 ones[2] VGND 0.769988f
C2110 rst VGND 0.724657f
C2111 pulse VGND 0.674805f
C2112 ones[7] VGND 0.486594f
C2113 ready VGND 0.568889f
C2114 ones[6] VGND 1.36849f
C2115 clk VGND 2.27788f
C2116 ones[3] VGND 0.389191f
C2117 ones[1] VGND 0.471797f
C2118 ones[8] VGND 0.452614f
C2119 ones[5] VGND 0.513732f
C2120 ones[0] VGND 0.798767f
C2121 ones[4] VGND 0.436512f
C2122 ones[9] VGND 0.731884f
C2123 ones[10] VGND 0.681711f
C2124 VPWR VGND 0.325241p
C2125 a_10199_2197# VGND 0.363289f
C2126 a_9871_2223# VGND 0.243145f
C2127 a_7123_2223# VGND 0.276055f
C2128 a_7194_2197# VGND 0.232044f
C2129 a_6987_2197# VGND 0.535606f
C2130 a_6994_2497# VGND 0.394413f
C2131 a_6703_2197# VGND 0.286403f
C2132 a_6607_2375# VGND 0.39011f
C2133 a_4363_2223# VGND 0.259894f
C2134 a_4434_2197# VGND 0.210268f
C2135 a_4227_2197# VGND 0.523746f
C2136 a_4234_2497# VGND 0.318743f
C2137 a_3943_2197# VGND 0.277976f
C2138 a_3847_2375# VGND 0.3671f
C2139 a_3187_2251# VGND 0.266352f
C2140 a_10039_3087# VGND 0.281338f
C2141 a_9595_3087# VGND 0.302276f
C2142 a_8907_2986# VGND 0.234704f
C2143 a_8631_2986# VGND 0.224914f
C2144 a_7847_3133# VGND 0.279117f
C2145 a_5363_2880# VGND 0.268162f
C2146 _065_ VGND 0.380497f
C2147 a_4771_2741# VGND 0.237535f
C2148 a_4111_2767# VGND 0.258427f
C2149 a_4279_2741# VGND 0.329287f
C2150 a_3686_2767# VGND 0.198071f
C2151 a_3854_2741# VGND 0.239878f
C2152 a_3413_2773# VGND 0.31047f
C2153 _014_ VGND 0.467812f
C2154 a_3247_2773# VGND 0.461894f
C2155 a_2866_3087# VGND 0.276258f
C2156 a_8076_3311# VGND 0.22038f
C2157 a_10199_3285# VGND 0.35399f
C2158 a_9921_3476# VGND 0.233105f
C2159 a_9213_3463# VGND 0.224859f
C2160 a_7886_3311# VGND 0.255271f
C2161 a_6871_3677# VGND 0.25302f
C2162 a_7039_3579# VGND 0.331714f
C2163 a_6446_3677# VGND 0.204369f
C2164 a_6614_3423# VGND 0.242953f
C2165 a_6173_3311# VGND 0.317034f
C2166 a_6007_3311# VGND 0.476503f
C2167 a_5399_3677# VGND 0.271521f
C2168 a_5567_3579# VGND 0.347859f
C2169 a_4974_3677# VGND 0.207244f
C2170 a_5142_3423# VGND 0.256736f
C2171 a_4701_3311# VGND 0.307329f
C2172 a_4535_3311# VGND 0.503758f
C2173 a_2682_3311# VGND 0.29856f
C2174 _013_ VGND 1.15133f
C2175 a_9919_4087# VGND 0.26206f
C2176 a_9079_3855# VGND 0.259518f
C2177 a_9247_3829# VGND 0.351699f
C2178 a_8654_3855# VGND 0.202571f
C2179 a_8822_3829# VGND 0.248608f
C2180 a_8381_3861# VGND 0.3067f
C2181 _015_ VGND 0.475863f
C2182 a_8215_3861# VGND 0.476511f
C2183 a_7847_3855# VGND 0.253792f
C2184 a_7111_4221# VGND 0.362977f
C2185 a_6515_4074# VGND 0.263866f
C2186 a_5717_4087# VGND 0.219855f
C2187 a_4731_4233# VGND 0.242088f
C2188 a_4802_4132# VGND 0.198229f
C2189 a_4602_3977# VGND 0.30661f
C2190 a_4595_4073# VGND 0.459966f
C2191 a_4311_4087# VGND 0.272459f
C2192 a_4215_4087# VGND 0.365003f
C2193 a_2879_3855# VGND 0.235551f
C2194 a_2460_3971# VGND 0.226241f
C2195 a_10147_4399# VGND 0.230341f
C2196 a_9687_4399# VGND 0.247017f
C2197 a_9096_4373# VGND 0.320688f
C2198 a_8459_4551# VGND 0.262634f
C2199 a_7980_4649# VGND 0.217269f
C2200 a_7239_4765# VGND 0.263404f
C2201 a_7407_4667# VGND 0.44336f
C2202 a_6814_4765# VGND 0.202208f
C2203 a_6982_4511# VGND 0.252315f
C2204 a_6541_4399# VGND 0.319426f
C2205 a_6375_4399# VGND 0.512767f
C2206 a_5675_4765# VGND 0.268436f
C2207 a_5843_4667# VGND 0.433273f
C2208 a_5250_4765# VGND 0.195245f
C2209 a_5418_4511# VGND 0.243927f
C2210 a_4977_4399# VGND 0.304756f
C2211 a_4811_4399# VGND 0.490928f
C2212 _076_ VGND 1.88245f
C2213 a_2509_4663# VGND 0.264169f
C2214 a_2409_4445# VGND 0.201544f
C2215 a_1867_4399# VGND 0.253866f
C2216 a_9815_4943# VGND 0.259503f
C2217 a_9983_4917# VGND 0.347788f
C2218 a_9390_4943# VGND 0.195572f
C2219 a_9558_4917# VGND 0.240008f
C2220 a_9117_4949# VGND 0.298816f
C2221 _016_ VGND 0.357967f
C2222 a_8951_4949# VGND 0.4642f
C2223 _046_ VGND 0.286721f
C2224 a_8447_5175# VGND 0.244437f
C2225 a_7419_5281# VGND 0.267031f
C2226 a_5960_5175# VGND 0.204882f
C2227 _075_ VGND 0.586587f
C2228 _085_ VGND 1.12082f
C2229 a_5687_5175# VGND 0.224201f
C2230 a_5141_4917# VGND 0.266393f
C2231 a_4627_5056# VGND 0.232375f
C2232 _083_ VGND 0.730277f
C2233 a_3983_5056# VGND 0.251415f
C2234 _063_ VGND 1.72951f
C2235 _062_ VGND 3.41367f
C2236 a_3611_4943# VGND 0.216177f
C2237 a_3431_4943# VGND 0.235939f
C2238 a_2823_4943# VGND 0.284028f
C2239 a_2991_4917# VGND 0.361021f
C2240 a_2398_4943# VGND 0.19621f
C2241 a_2566_4917# VGND 0.252225f
C2242 a_2125_4949# VGND 0.326793f
C2243 a_1959_4949# VGND 0.459042f
C2244 a_1499_5056# VGND 0.238262f
C2245 net11 VGND 3.17809f
C2246 a_9515_5487# VGND 0.244644f
C2247 a_9586_5461# VGND 0.200962f
C2248 a_9379_5461# VGND 0.491437f
C2249 a_9386_5761# VGND 0.298603f
C2250 a_9095_5461# VGND 0.263434f
C2251 a_8999_5639# VGND 0.3486f
C2252 a_8109_5639# VGND 0.229851f
C2253 a_7331_5853# VGND 0.262513f
C2254 a_7499_5755# VGND 0.459311f
C2255 a_6906_5853# VGND 0.192291f
C2256 a_7074_5599# VGND 0.244139f
C2257 a_6633_5487# VGND 0.306038f
C2258 a_6467_5487# VGND 0.475482f
C2259 a_4697_5461# VGND 2.03774f
C2260 _000_ VGND 0.497359f
C2261 _082_ VGND 0.885901f
C2262 a_10287_6250# VGND 0.239222f
C2263 a_9915_6337# VGND 0.229064f
C2264 a_9739_6005# VGND 0.211519f
C2265 a_8779_6409# VGND 0.241103f
C2266 a_8850_6308# VGND 0.20255f
C2267 a_8650_6153# VGND 0.311672f
C2268 a_8643_6249# VGND 0.456654f
C2269 a_8359_6263# VGND 0.260803f
C2270 a_8263_6263# VGND 0.352072f
C2271 a_7939_6031# VGND 0.245314f
C2272 a_7239_6031# VGND 0.273421f
C2273 a_7407_6005# VGND 0.454697f
C2274 a_6814_6031# VGND 0.196413f
C2275 a_6982_6005# VGND 0.250201f
C2276 a_6541_6037# VGND 0.355561f
C2277 a_6375_6037# VGND 0.491132f
C2278 a_4627_6031# VGND 0.242435f
C2279 _061_ VGND 0.320809f
C2280 _091_ VGND 0.942162f
C2281 a_3797_6147# VGND 0.242372f
C2282 _081_ VGND 0.559394f
C2283 a_3697_6031# VGND 0.205147f
C2284 _049_ VGND 1.90307f
C2285 a_3029_6031# VGND 0.359747f
C2286 a_1670_6351# VGND 0.299695f
C2287 counter\[7\] VGND 1.72316f
C2288 _007_ VGND 0.861672f
C2289 a_9515_6575# VGND 0.240214f
C2290 a_9586_6549# VGND 0.196227f
C2291 a_9379_6549# VGND 0.483223f
C2292 a_9386_6849# VGND 0.300555f
C2293 a_9095_6549# VGND 0.255934f
C2294 a_8999_6727# VGND 0.339398f
C2295 a_8175_6549# VGND 0.256461f
C2296 a_6169_6549# VGND 1.99459f
C2297 a_5087_6575# VGND 0.238726f
C2298 _054_ VGND 0.353882f
C2299 _058_ VGND 1.2044f
C2300 a_2247_6575# VGND 0.241305f
C2301 a_2318_6549# VGND 0.204031f
C2302 a_2111_6549# VGND 0.511761f
C2303 a_2118_6849# VGND 0.315704f
C2304 a_1827_6549# VGND 0.26767f
C2305 a_1731_6727# VGND 0.350803f
C2306 _020_ VGND 1.3302f
C2307 a_5261_7439# VGND 0.188513f
C2308 _043_ VGND 3.10846f
C2309 _051_ VGND 0.343788f
C2310 a_10195_7338# VGND 0.23819f
C2311 a_8390_7119# VGND 1.90006f
C2312 clknet_0_clk VGND 2.52641f
C2313 a_7663_7485# VGND 0.273016f
C2314 _024_ VGND 1.06466f
C2315 a_4535_7232# VGND 0.237639f
C2316 a_4073_7235# VGND 0.249223f
C2317 _044_ VGND 0.800827f
C2318 a_3973_7119# VGND 0.216662f
C2319 net10 VGND 1.37606f
C2320 a_2639_7119# VGND 0.289445f
C2321 a_2807_7093# VGND 0.361582f
C2322 a_2214_7119# VGND 0.199234f
C2323 a_2382_7093# VGND 0.259329f
C2324 a_1941_7125# VGND 0.331668f
C2325 a_1775_7125# VGND 0.516235f
C2326 _038_ VGND 0.738197f
C2327 a_6283_7669# VGND 0.284426f
C2328 _011_ VGND 0.831904f
C2329 counter\[6\] VGND 3.05582f
C2330 _074_ VGND 2.05815f
C2331 _037_ VGND 4.39241f
C2332 a_10239_7663# VGND 0.221651f
C2333 a_9963_7663# VGND 0.209472f
C2334 a_9687_7663# VGND 0.244029f
C2335 a_6475_7913# VGND 0.255617f
C2336 _093_ VGND 1.97153f
C2337 _092_ VGND 0.350828f
C2338 a_4668_7913# VGND 0.227025f
C2339 a_1991_7691# VGND 0.280914f
C2340 _069_ VGND 0.641685f
C2341 _004_ VGND 0.514413f
C2342 a_9832_8181# VGND 0.333603f
C2343 a_9503_8207# VGND 0.215976f
C2344 _077_ VGND 0.833746f
C2345 _078_ VGND 1.78926f
C2346 a_9091_8439# VGND 0.240883f
C2347 a_8720_8439# VGND 0.204585f
C2348 _027_ VGND 1.17165f
C2349 _029_ VGND 0.695902f
C2350 _019_ VGND 0.425257f
C2351 _033_ VGND 1.51317f
C2352 a_8447_8439# VGND 0.244365f
C2353 a_6007_8207# VGND 0.257044f
C2354 _048_ VGND 0.696553f
C2355 a_4580_8439# VGND 0.209537f
C2356 _035_ VGND 0.655076f
C2357 _036_ VGND 0.687851f
C2358 _021_ VGND 0.849366f
C2359 a_4307_8439# VGND 0.244029f
C2360 _053_ VGND 1.49089f
C2361 _052_ VGND 4.52867f
C2362 _050_ VGND 5.84785f
C2363 a_9624_8751# VGND 0.165974f
C2364 a_9533_8751# VGND 0.128869f
C2365 _010_ VGND 0.77489f
C2366 _006_ VGND 2.03472f
C2367 a_10239_8751# VGND 0.238834f
C2368 net9 VGND 1.88835f
C2369 a_9435_9001# VGND 0.233283f
C2370 _079_ VGND 0.468812f
C2371 a_8447_8916# VGND 0.24948f
C2372 a_7699_9117# VGND 0.28692f
C2373 a_7867_9019# VGND 0.453022f
C2374 a_7274_9117# VGND 0.203681f
C2375 a_7442_8863# VGND 0.277015f
C2376 a_7001_8751# VGND 0.327182f
C2377 _022_ VGND 0.76076f
C2378 a_6835_8751# VGND 0.487851f
C2379 net2 VGND 2.1247f
C2380 _025_ VGND 2.631f
C2381 a_4120_8731# VGND 0.206268f
C2382 _088_ VGND 0.983637f
C2383 a_4521_8903# VGND 0.242711f
C2384 _087_ VGND 1.10502f
C2385 _026_ VGND 4.01319f
C2386 _017_ VGND 0.684376f
C2387 a_3847_8903# VGND 0.250049f
C2388 a_2971_8751# VGND 0.405212f
C2389 _039_ VGND 3.3036f
C2390 _041_ VGND 1.85666f
C2391 _001_ VGND 0.705171f
C2392 _009_ VGND 1.10282f
C2393 a_7791_9295# VGND 0.26301f
C2394 a_7959_9269# VGND 0.351514f
C2395 a_7366_9295# VGND 0.208052f
C2396 a_7534_9269# VGND 0.260917f
C2397 a_7093_9301# VGND 0.330431f
C2398 _012_ VGND 0.691647f
C2399 a_6927_9301# VGND 0.513621f
C2400 a_4903_9295# VGND 0.28119f
C2401 _064_ VGND 0.643357f
C2402 _089_ VGND 0.359705f
C2403 a_4123_9514# VGND 0.261802f
C2404 _059_ VGND 2.24176f
C2405 a_1460_9269# VGND 0.39426f
C2406 a_10239_9839# VGND 0.240725f
C2407 _067_ VGND 7.70081f
C2408 a_9091_10004# VGND 0.271773f
C2409 _066_ VGND 1.06953f
C2410 _090_ VGND 0.857707f
C2411 net1 VGND 4.10642f
C2412 net14 VGND 3.30797f
C2413 _023_ VGND 1.86112f
C2414 _047_ VGND 2.85162f
C2415 _008_ VGND 2.17184f
C2416 a_6939_9839# VGND 0.241971f
C2417 a_7010_9813# VGND 0.198677f
C2418 a_6803_9813# VGND 0.513919f
C2419 a_6810_10113# VGND 0.311987f
C2420 a_6519_9813# VGND 0.25673f
C2421 a_6423_9991# VGND 0.349961f
C2422 a_5785_9813# VGND 0.270868f
C2423 a_4981_9991# VGND 0.238563f
C2424 _042_ VGND 2.78071f
C2425 _040_ VGND 0.947272f
C2426 net12 VGND 2.61782f
C2427 a_1461_9813# VGND 0.286092f
C2428 _032_ VGND 0.818694f
C2429 _018_ VGND 1.87403f
C2430 _034_ VGND 1.61808f
C2431 counter\[5\] VGND 1.72876f
C2432 _056_ VGND 0.733902f
C2433 _086_ VGND 1.96464f
C2434 a_10239_10383# VGND 0.244022f
C2435 net8 VGND 4.39882f
C2436 a_8215_10496# VGND 0.2557f
C2437 _031_ VGND 1.93035f
C2438 _030_ VGND 0.573043f
C2439 _028_ VGND 5.30797f
C2440 clknet_1_1__leaf_clk VGND 3.68688f
C2441 _002_ VGND 0.336239f
C2442 a_7307_10761# VGND 0.239014f
C2443 a_7378_10660# VGND 0.201799f
C2444 a_7178_10505# VGND 0.322248f
C2445 a_7171_10601# VGND 0.489319f
C2446 a_6887_10615# VGND 0.250305f
C2447 a_6719_10615# VGND 0.419081f
C2448 _045_ VGND 0.565812f
C2449 a_6425_10602# VGND 0.22725f
C2450 net7 VGND 3.25618f
C2451 net6 VGND 5.70483f
C2452 net5 VGND 2.99093f
C2453 net3 VGND 5.55466f
C2454 a_5507_10357# VGND 0.253769f
C2455 clknet_1_0__leaf_clk VGND 4.84413f
C2456 _005_ VGND 2.29516f
C2457 a_3811_10761# VGND 0.254111f
C2458 a_3882_10660# VGND 0.217938f
C2459 a_3682_10505# VGND 0.326128f
C2460 a_3675_10601# VGND 0.528106f
C2461 a_3391_10615# VGND 0.269835f
C2462 a_3295_10615# VGND 0.360812f
C2463 counter\[0\] VGND 3.7463f
C2464 a_2555_10704# VGND 0.323382f
C2465 counter\[3\] VGND 3.03877f
C2466 counter\[2\] VGND 7.15489f
C2467 counter\[1\] VGND 3.91861f
C2468 a_2191_10615# VGND 0.206505f
C2469 a_1683_10496# VGND 0.255933f
C2470 _055_ VGND 1.65521f
C2471 _084_ VGND 2.06894f
C2472 counter\[4\] VGND 5.4164f
C2473 _068_ VGND 5.30438f
C2474 counter\[9\] VGND 5.48646f
C2475 counter\[10\] VGND 1.99113f
C2476 _057_ VGND 5.34439f
C2477 _073_ VGND 1.15186f
C2478 _072_ VGND 0.996701f
C2479 _060_ VGND 3.96885f
C2480 _071_ VGND 1.92234f
C2481 _003_ VGND 2.32735f
C2482 a_10239_10927# VGND 0.260755f
C2483 net13 VGND 5.60681f
C2484 _080_ VGND 6.04496f
C2485 counter\[8\] VGND 3.97778f
C2486 a_9687_10927# VGND 0.25606f
C2487 net4 VGND 3.54498f
C2488 a_8256_11177# VGND 0.248046f
C2489 a_6423_11079# VGND 0.286402f
C2490 a_3799_10927# VGND 0.273406f
C2491 a_2603_10927# VGND 0.29171f
C2492 _070_ VGND 2.15177f
.ends

