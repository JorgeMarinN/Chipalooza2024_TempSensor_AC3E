magic
tech sky130A
magscale 1 2
timestamp 1713593032
<< error_p >>
rect -29 -107 29 -101
rect -29 -141 -17 -107
rect -29 -147 29 -141
<< pwell >>
rect -99 -95 99 157
<< nmos >>
rect -15 -69 15 131
<< ndiff >>
rect -73 116 -15 131
rect -73 82 -61 116
rect -27 82 -15 116
rect -73 48 -15 82
rect -73 14 -61 48
rect -27 14 -15 48
rect -73 -20 -15 14
rect -73 -54 -61 -20
rect -27 -54 -15 -20
rect -73 -69 -15 -54
rect 15 116 73 131
rect 15 82 27 116
rect 61 82 73 116
rect 15 48 73 82
rect 15 14 27 48
rect 61 14 73 48
rect 15 -20 73 14
rect 15 -54 27 -20
rect 61 -54 73 -20
rect 15 -69 73 -54
<< ndiffc >>
rect -61 82 -27 116
rect -61 14 -27 48
rect -61 -54 -27 -20
rect 27 82 61 116
rect 27 14 61 48
rect 27 -54 61 -20
<< poly >>
rect -15 131 15 157
rect -15 -91 15 -69
rect -33 -107 33 -91
rect -33 -141 -17 -107
rect 17 -141 33 -107
rect -33 -157 33 -141
<< polycont >>
rect -17 -141 17 -107
<< locali >>
rect -61 116 -27 135
rect -61 48 -27 50
rect -61 12 -27 14
rect -61 -73 -27 -54
rect 27 116 61 135
rect 27 48 61 50
rect 27 12 61 14
rect 27 -73 61 -54
rect -33 -141 -17 -107
rect 17 -141 33 -107
<< viali >>
rect -61 82 -27 84
rect -61 50 -27 82
rect -61 -20 -27 12
rect -61 -22 -27 -20
rect 27 82 61 84
rect 27 50 61 82
rect 27 -20 61 12
rect 27 -22 61 -20
rect -17 -141 17 -107
<< metal1 >>
rect -67 84 -21 131
rect -67 50 -61 84
rect -27 50 -21 84
rect -67 12 -21 50
rect -67 -22 -61 12
rect -27 -22 -21 12
rect -67 -69 -21 -22
rect 21 84 67 131
rect 21 50 27 84
rect 61 50 67 84
rect 21 12 67 50
rect 21 -22 27 12
rect 61 -22 67 12
rect 21 -69 67 -22
rect -29 -107 29 -101
rect -29 -141 -17 -107
rect 17 -141 29 -107
rect -29 -147 29 -141
<< end >>
