* NGSPICE file created from ONES_COUNTER_pex.ext - technology: sky130A

.subckt ONES_COUNTER_pex VGND VPWR clk rst pulse ready ones[0] ones[1] ones[2] ones[3] ones[4] ones[5]
+ ones[6] ones[7] ones[8] ones[9] ones[10]
X0 a_2957_2999# counter\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X1 a_1832_6825# counter\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.33 w=0.42 l=0.15
X2 VPWR _033_ a_8352_9527# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X3 a_9183_8573# a_8963_8585# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.08 w=0.42 l=0.15
X4 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=135 ps=1.29k w=0.87 l=0.59
X5 VPWR net14 a_9810_6147# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.33 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 a_3368_6351# _087_ a_3277_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0991 ps=0.955 w=0.65 l=0.15
X7 a_6546_5487# net8 a_6377_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X8 VGND a_5383_2741# a_5341_3145# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X9 a_9305_10927# _019_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X10 a_6701_6369# net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X11 a_2879_9839# net5 a_2773_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X12 VGND a_1669_6727# _083_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X13 a_8942_5220# a_8735_5161# a_9118_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0766 ps=0.785 w=0.42 l=0.15
X14 VGND clknet_1_1__leaf_clk a_8951_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X15 a_9919_8439# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X16 _059_ net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VPWR _031_ a_2877_4649# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 clknet_1_1__leaf_clk a_8022_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 VGND a_9558_11039# a_9516_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0696 ps=0.765 w=0.42 l=0.15
X20 _030_ a_2736_5059# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X21 ones[10] a_8307_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X22 a_2691_6825# _043_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X23 VGND a_3330_7396# a_3259_7497# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0989 ps=0.995 w=0.64 l=0.15
X24 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X25 a_9919_8439# _060_ a_10153_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X26 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=86.8 ps=916 w=0.55 l=0.59
X27 a_8022_7119# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X28 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X29 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X30 VPWR clknet_1_1__leaf_clk a_6007_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X31 a_8815_9527# a_9088_9527# a_9046_9655# VGND sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X32 VPWR _043_ a_7111_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X33 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X34 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X35 VPWR a_5326_7093# a_5253_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0766 ps=0.785 w=0.42 l=0.15
X36 VGND a_9827_7351# _082_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X37 VPWR clknet_1_1__leaf_clk a_8951_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X38 a_1761_2767# _007_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X39 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X40 VPWR pulse a_1407_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.32 as=0.265 ps=2.53 w=1 l=0.15
X41 VPWR _001_ a_2481_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X42 VGND counter\[3\] a_2472_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X43 a_4169_9001# counter\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X44 a_1925_2473# net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X45 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X46 VPWR a_6527_6263# _042_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X47 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X48 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X49 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X50 VGND a_4227_5161# a_4234_5065# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X51 a_5253_7119# a_4719_7125# a_5158_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.0682 ps=0.745 w=0.42 l=0.15
X52 a_4319_7637# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X53 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X54 _074_ a_5915_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.33 w=1 l=0.15
X55 a_2849_6397# _065_ a_2777_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X56 VPWR a_4227_9513# a_4234_9417# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X57 clknet_1_0__leaf_clk a_4053_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X58 VPWR a_7258_4511# a_7185_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0766 ps=0.785 w=0.42 l=0.15
X59 a_4434_5220# a_4227_5161# a_4610_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0766 ps=0.785 w=0.42 l=0.15
X60 a_3481_9867# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X61 ones[8] a_9963_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X62 VGND _004_ a_4873_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X63 _052_ net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X64 a_6503_3677# a_5639_3311# a_6246_3423# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.07 w=0.42 l=0.15
X65 a_7469_10703# net4 a_7385_10703# VGND sky130_fd_pr__nfet_01v8 ad=0.184 pd=1.21 as=0.0877 ps=0.92 w=0.65 l=0.15
X66 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X67 VPWR net9 a_3215_4551# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X68 counter\[7\] a_2439_2741# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X69 a_5941_5309# _037_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X70 VPWR a_7895_8916# _008_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X71 _017_ _041_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X72 _061_ a_3243_11293# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.228 ps=1.74 w=1 l=0.15
X73 VGND net4 a_8307_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X74 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X75 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X76 a_7185_4765# a_6651_4399# a_7090_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.0682 ps=0.745 w=0.42 l=0.15
X77 a_4610_4943# a_4363_5321# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X78 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X79 VGND _043_ a_5537_5263# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X80 a_6069_5487# counter\[4\] a_5997_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X81 a_8942_5220# a_8742_5065# a_9091_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X82 a_4322_10927# counter\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.175 ps=1.26 w=0.42 l=0.15
X83 counter\[2\] a_8143_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X84 a_7975_6031# a_7111_6037# a_7718_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.07 w=0.42 l=0.15
X85 VPWR _060_ a_9827_7351# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X86 a_7550_6031# a_7111_6037# a_7465_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X87 VPWR counter\[3\] a_1665_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.128 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X88 a_6835_3968# _083_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X89 a_8355_5175# a_8451_5175# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X90 clknet_1_1__leaf_clk a_8022_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X91 _056_ a_1665_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.103 ps=1 w=0.65 l=0.15
X92 a_2589_4221# net7 a_2501_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X93 _085_ a_6835_3968# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.33 w=1 l=0.15
X94 a_4958_2741# a_4790_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.08 w=0.64 l=0.15
X95 a_1573_8213# a_1407_8213# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X96 ones[6] a_10239_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X97 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X98 ones[2] a_10239_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X99 VGND _059_ a_6375_2775# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X100 VGND _078_ a_5057_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X101 VPWR a_4053_6005# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X102 VGND a_6607_5175# counter\[10\] VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X103 a_1748_5303# _069_ a_1676_5303# VGND sky130_fd_pr__nfet_01v8 ad=0.0535 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X104 VPWR a_2134_5461# a_2063_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.07 w=0.75 l=0.15
X105 a_4781_6575# a_4234_6849# a_4434_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0682 ps=0.745 w=0.42 l=0.15
X106 a_4162_6575# a_3847_6727# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X107 VGND a_2473_6549# _049_ VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X108 VPWR a_6671_3579# a_6587_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X109 VGND a_3847_6727# counter\[3\] VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X110 a_4675_7663# a_4455_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.08 w=0.42 l=0.15
X111 VGND _050_ a_4505_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X112 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X113 VPWR _026_ _031_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X114 a_7676_6409# a_7277_6037# a_7550_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X115 a_3220_9655# _027_ a_3148_9655# VGND sky130_fd_pr__nfet_01v8 ad=0.0535 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X116 VGND counter\[1\] a_1941_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.103 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X117 a_5411_7815# a_5684_7643# a_5642_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X118 VGND a_7895_8916# _008_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X119 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X120 a_3943_5175# a_4234_5065# a_4185_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X121 VPWR counter\[9\] a_5607_11079# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X122 a_7123_5321# a_6987_5161# a_6703_5175# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
X123 a_9558_11039# a_9390_11293# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.08 w=0.64 l=0.15
X124 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X125 VPWR a_8942_5220# a_8871_5321# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.07 w=0.75 l=0.15
X126 VGND clknet_1_1__leaf_clk a_6559_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X128 net5 a_2439_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X129 a_10245_5309# _030_ a_10173_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X130 a_9135_5737# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.148 ps=1.29 w=1 l=0.15
X131 _067_ a_2695_6144# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X132 a_4526_7637# a_4326_7937# a_4675_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X133 a_4434_5220# a_4234_5065# a_4583_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X134 VPWR counter\[0\] a_9137_7913# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X135 _012_ _025_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.0877 ps=0.92 w=0.65 l=0.15
X136 a_3259_7497# a_3123_7337# a_2839_7351# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
X137 a_6817_4399# a_6651_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X138 a_3775_9527# a_3943_9527# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X139 a_5993_3311# _016_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X140 a_5215_2767# a_4351_2773# a_4958_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.07 w=0.42 l=0.15
X141 a_3847_5175# a_3943_5175# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X142 clknet_1_0__leaf_clk a_4053_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X143 _072_ a_1632_3971# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X145 clknet_0_clk a_5722_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X146 VPWR clknet_1_0__leaf_clk a_5639_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X147 VGND a_4434_5220# a_4363_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0989 ps=0.995 w=0.64 l=0.15
X148 a_9275_6263# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.33 w=0.42 l=0.15
X149 a_4873_7663# a_4319_7637# a_4526_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X150 a_4781_5321# a_4227_5161# a_4434_5220# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X151 clknet_1_0__leaf_clk a_4053_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X152 VGND a_8022_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X153 a_4790_2767# a_4351_2773# a_4705_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X154 VGND counter\[5\] a_4338_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X155 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X156 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X157 _062_ counter\[1\] a_1861_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X158 VPWR clknet_1_0__leaf_clk a_1407_8213# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X159 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X160 a_1632_3971# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X161 VPWR a_2439_2741# a_2355_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X162 _050_ net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.215 ps=1.43 w=1 l=0.15
X163 VPWR a_7255_3285# _054_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X164 _012_ _025_ a_9411_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X165 clknet_0_clk a_5722_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X166 VGND a_6987_5161# a_6994_5065# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X167 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X168 VPWR a_1547_10004# _007_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X169 net7 a_7039_9019# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X170 a_4916_3145# a_4517_2773# a_4790_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X171 VPWR _028_ a_4627_8320# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X172 a_1547_10004# _082_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X173 a_9209_10389# a_9043_10389# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X174 clknet_1_1__leaf_clk a_8022_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X175 a_6871_9117# a_6173_8751# a_6614_8863# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X176 VPWR _055_ a_3307_9991# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X177 VGND clknet_1_0__leaf_clk a_1407_2773# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X178 VPWR a_5383_2741# a_5299_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X179 a_5709_7497# a_4719_7125# a_5583_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X180 VPWR a_3939_7815# counter\[4\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X181 VPWR net14 _091_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X182 a_4709_8573# _028_ a_4627_8320# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X183 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X184 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X185 VGND a_4053_6005# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X186 VGND _080_ a_1669_6727# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X187 VPWR a_3330_7396# a_3259_7497# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.07 w=0.75 l=0.15
X188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X189 ones[8] a_9963_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X190 a_7951_5487# a_7822_5761# a_7531_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X191 a_7531_5461# a_7822_5761# a_7773_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X192 VPWR a_2014_8181# a_1941_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0766 ps=0.785 w=0.42 l=0.15
X193 _091_ net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X194 VGND a_1407_10927# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X195 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X196 a_8009_3145# a_7019_2773# a_7883_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X197 VPWR _030_ a_10011_5175# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X198 a_5215_2767# a_4517_2773# a_4958_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X199 VPWR _021_ a_9289_5321# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X200 a_8963_8585# a_8834_8329# a_8543_8439# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X201 a_7373_2767# _015_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X202 VGND a_8051_2741# a_8009_3145# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X203 VPWR counter\[1\] _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X204 _026_ a_9655_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X205 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X206 a_3058_7485# a_2743_7351# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X207 a_1643_5461# a_1927_5461# a_1862_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X208 VGND a_6803_9513# a_6810_9417# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X209 VPWR net13 a_8583_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X210 VPWR a_8079_5162# _004_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X211 VPWR counter\[3\] a_4043_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X212 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X213 VGND a_5722_6575# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X214 a_7185_2773# a_7019_2773# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X215 VPWR a_7815_5461# a_7822_5761# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X216 a_2736_9001# _039_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X217 clknet_1_0__leaf_clk a_4053_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X218 a_9279_8725# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X219 net7 a_7039_9019# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X220 _031_ net7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X221 _015_ a_2971_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X222 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X223 ones[6] a_10239_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X224 a_8369_5487# a_7815_5461# a_8022_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X226 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X227 a_6423_9527# a_6519_9527# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X228 a_7255_3285# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.228 ps=1.74 w=0.42 l=0.15
X229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X230 a_2115_2223# net3 a_1925_2473# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X231 VPWR _009_ a_4781_5321# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X232 _068_ a_4043_10901# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X233 _038_ a_2795_4649# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X234 a_4455_7663# a_4326_7937# a_4035_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X235 a_4363_5321# a_4234_5065# a_3943_5175# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X236 a_5779_5175# _023_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X237 VGND a_3939_7815# counter\[4\] VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X238 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X240 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X241 clknet_1_1__leaf_clk a_8022_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X242 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X243 _021_ _053_ a_9135_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X244 a_4434_9572# a_4234_9417# a_4583_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X245 clknet_1_1__leaf_clk a_8022_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X246 a_3123_7337# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X247 a_9034_8484# a_8827_8425# a_9210_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0766 ps=0.785 w=0.42 l=0.15
X248 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X249 a_1489_4943# _068_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X250 VPWR a_7363_5461# counter\[0\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X251 VPWR a_7619_8916# _009_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X252 net3 a_3775_9527# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X253 VGND net13 a_8583_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X254 a_9558_11039# a_9390_11293# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.179 ps=1.26 w=0.75 l=0.15
X255 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X256 a_9571_8751# _037_ a_9475_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X257 a_6361_8751# _014_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X258 VPWR a_2472_10901# _069_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X259 a_6089_9615# counter\[4\] _071_ VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X260 VPWR a_6607_5175# counter\[10\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X261 VGND a_1927_5461# a_1934_5761# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X262 a_4035_7637# a_4326_7937# a_4277_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X263 VGND a_9034_8484# a_8963_8585# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0989 ps=0.995 w=0.64 l=0.15
X264 net5 a_2439_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X265 _011_ _093_ a_4909_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X266 _070_ a_1589_5059# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.33 w=1 l=0.15
X267 a_4434_9572# a_4227_9513# a_4610_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0766 ps=0.785 w=0.42 l=0.15
X268 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X269 _062_ counter\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X270 a_6446_9117# a_6007_8751# a_6361_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X271 VGND a_4053_6005# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X272 VPWR a_5722_6575# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X273 a_9210_8207# a_8963_8585# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X274 VGND counter\[6\] a_9544_3561# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X275 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X276 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X277 a_2818_5059# _026_ a_2736_5059# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X278 _016_ a_5126_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X279 a_4227_6549# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X280 a_4781_9673# a_4227_9513# a_4434_9572# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X281 VGND _028_ a_3220_9655# VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0535 ps=0.675 w=0.42 l=0.15
X282 VGND _080_ a_10100_7351# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X283 VPWR a_2743_7351# net6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X284 a_5216_5487# _028_ a_5126_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.114 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X285 net13 a_10075_10357# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X286 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X287 _005_ a_6375_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X288 a_8198_5853# a_7951_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X289 _047_ a_3970_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X290 _022_ a_1867_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X291 a_4610_9295# a_4363_9673# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X293 VPWR net11 _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.215 pd=1.43 as=0.135 ps=1.27 w=1 l=0.15
X294 VGND _024_ _012_ VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.17 w=0.65 l=0.15
X295 a_1885_5853# a_1475_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X296 VGND counter\[2\] a_6093_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X297 VGND clknet_0_clk a_8022_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X298 a_6572_8751# a_6173_8751# a_6446_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X299 a_5264_2229# a_5077_2269# a_5177_2487# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X300 a_7549_9839# a_6559_9839# a_7423_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X301 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X302 a_9437_6397# _026_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X303 a_6519_9527# a_6810_9417# a_6761_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X304 VGND a_5722_6575# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X305 a_4227_5161# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X306 _079_ a_4903_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X307 VGND a_10075_10357# a_10033_10761# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X308 a_9711_2767# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X309 VGND _074_ a_5684_7643# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X310 VPWR net8 a_10239_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X311 _055_ a_8583_6397# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X312 VPWR a_8022_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X313 clknet_1_0__leaf_clk a_4053_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X314 a_4985_4399# _060_ a_4903_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X315 VGND a_7619_8916# _009_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X316 VGND a_8022_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0578 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X317 a_8965_9655# _044_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0535 pd=0.675 as=0.122 ps=1.08 w=0.42 l=0.15
X318 VPWR a_7883_2767# a_8051_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X319 VGND rst a_1407_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0682 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X320 net9 a_6671_3579# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X321 a_8859_6397# counter\[7\] a_8753_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X322 VGND a_6614_8863# a_6572_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0696 ps=0.765 w=0.42 l=0.15
X323 VPWR _067_ a_6099_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X324 VPWR _078_ a_4903_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X325 VGND _037_ a_2603_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.157 pd=1.17 as=0.109 ps=1.36 w=0.42 l=0.15
X326 a_2537_10749# _072_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X327 a_3243_11293# a_3063_11293# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X328 VPWR net7 a_10239_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X329 a_7458_2767# a_7185_2773# a_7373_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X330 a_8369_5487# a_7822_5761# a_8022_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0682 ps=0.745 w=0.42 l=0.15
X331 a_3943_9527# a_4234_9417# a_4185_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X332 VPWR _055_ a_7527_4087# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X333 VGND a_7363_5461# counter\[0\] VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X334 a_6546_5487# _023_ a_6460_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X335 VPWR a_8263_6740# _003_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X336 VPWR counter\[1\] a_4043_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0745 ps=0.775 w=0.42 l=0.15
X337 a_4719_3311# _039_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X338 VGND a_8079_5162# _004_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X339 a_8447_8439# a_8543_8439# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X340 a_4227_6549# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X341 a_2397_8585# a_1407_8213# a_2271_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X342 clknet_1_1__leaf_clk a_8022_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X343 a_3277_6351# _060_ a_3179_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0991 pd=0.955 as=0.201 ps=1.92 w=0.65 l=0.15
X344 a_3120_2883# counter\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.146 ps=1.33 w=0.42 l=0.15
X345 VPWR _068_ a_4169_9001# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X346 a_5537_5263# net12 _046_ VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X347 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
D0 VGND net1 sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X348 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X349 VGND _003_ a_4781_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X350 a_3775_9527# a_3943_9527# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X351 a_3063_11293# counter\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X352 a_5993_3311# _016_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X353 _015_ a_2971_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X354 VGND a_7591_10107# a_7549_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X355 a_8355_5175# a_8451_5175# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X356 a_1927_5461# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X357 a_7010_9572# a_6810_9417# a_7159_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X358 a_2685_9839# net7 a_2603_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X359 a_6361_8751# _014_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X360 VPWR net13 _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0.135 ps=1.27 w=1 l=0.15
X361 VPWR clknet_1_1__leaf_clk a_6651_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X362 a_4162_5309# a_3847_5175# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X363 a_7541_5321# a_6994_5065# a_7194_5220# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0682 ps=0.745 w=0.42 l=0.15
X364 VPWR a_7626_2741# a_7553_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0766 ps=0.785 w=0.42 l=0.15
X365 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X366 VPWR a_8735_5161# a_8742_5065# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X367 a_7010_9572# a_6803_9513# a_7186_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0766 ps=0.785 w=0.42 l=0.15
X368 VPWR a_3123_7337# a_3130_7241# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X369 clknet_0_clk a_5722_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X370 a_4363_9673# a_4234_9417# a_3943_9527# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X371 VPWR net1 a_9711_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X372 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X373 a_7357_9673# a_6803_9513# a_7010_9572# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X374 _060_ a_6375_2775# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X375 _023_ a_3932_2883# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X376 a_2419_4221# net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X377 VGND a_5722_6575# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X378 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X379 VGND a_8815_9527# _045_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X380 a_7718_6005# a_7550_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.08 w=0.64 l=0.15
X381 VPWR a_9655_9813# _026_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.62 as=0.165 ps=1.33 w=1 l=0.15
X382 a_9711_2767# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X383 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X384 a_7553_2767# a_7019_2773# a_7458_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.0682 ps=0.745 w=0.42 l=0.15
X385 a_9306_7663# counter\[2\] a_9137_7913# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X386 a_7186_9295# a_6939_9673# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X387 VGND a_8022_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X389 a_6446_9117# a_6173_8751# a_6361_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X390 a_4583_6575# a_4363_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.08 w=0.42 l=0.15
X391 a_8815_9527# a_9088_9527# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X392 _010_ a_3179_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X393 a_1665_10383# counter\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.128 ps=1.03 w=0.42 l=0.15
X394 VPWR _088_ a_5177_2487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.0744 ps=0.815 w=0.42 l=0.15
X395 a_9126_3311# _023_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X396 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X397 a_1475_5461# a_1643_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X398 _028_ net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X399 _057_ a_3247_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X400 a_9650_10357# a_9482_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.179 ps=1.26 w=0.75 l=0.15
X401 a_9482_10383# a_9209_10389# a_9397_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X402 a_3847_5175# a_3943_5175# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X403 _065_ counter\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X404 _050_ net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X405 VPWR a_5383_2741# net14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X406 VPWR net11 a_2818_9001# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.33 as=0.0441 ps=0.63 w=0.42 l=0.15
X407 a_5781_10955# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X409 VPWR net5 a_9963_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X410 a_9589_6575# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X411 _063_ a_8624_10499# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.33 w=1 l=0.15
X412 VGND a_7010_9572# a_6939_9673# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0989 ps=0.995 w=0.64 l=0.15
X413 VGND a_9650_10357# a_9608_10761# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0696 ps=0.765 w=0.42 l=0.15
D1 VGND _086_ sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X414 a_4434_6549# a_4234_6849# a_4583_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X415 a_9907_10383# a_9209_10389# a_9650_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X416 VGND a_9275_6263# _033_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X417 _041_ _028_ a_2051_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X418 VPWR a_9919_8439# _064_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X419 VPWR clk a_5722_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X420 _022_ a_1867_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X421 a_4705_2767# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X422 a_8022_7119# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X423 net2 a_1407_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.32 w=1 l=0.15
X424 VPWR a_8079_9527# _036_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X425 VGND a_4864_3829# _027_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X426 VPWR clknet_1_0__leaf_clk a_4719_7125# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X427 a_6998_10205# a_6725_9839# a_6913_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X428 net11 a_7591_10107# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X429 a_8827_8425# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X430 a_7357_9673# a_6810_9417# a_7010_9572# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0682 ps=0.745 w=0.42 l=0.15
X431 _081_ a_6178_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X432 a_9043_3561# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.148 ps=1.29 w=1 l=0.15
X433 VPWR a_6614_8863# a_6541_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0766 ps=0.785 w=0.42 l=0.15
X434 VPWR net6 a_9655_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0745 ps=0.775 w=0.42 l=0.15
X435 VPWR net4 a_8307_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X436 VGND net8 a_10239_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X437 a_4781_6575# a_4227_6549# a_4434_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X438 VGND pulse a_1407_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0682 pd=0.745 as=0.111 ps=1.37 w=0.42 l=0.15
X439 VGND a_4053_6005# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X441 VPWR a_4043_10901# _068_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=1.62 as=0.165 ps=1.33 w=1 l=0.15
X442 VPWR _054_ a_1867_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X443 a_4517_2773# a_4351_2773# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X444 VPWR a_2439_8181# a_2355_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X445 VPWR _005_ a_9381_8585# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X446 VGND a_2375_10615# _073_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X447 a_7090_4765# a_6817_4399# a_7005_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X449 a_8693_4943# a_8355_5175# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X450 a_4524_10927# counter\[0\] a_4418_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.062 pd=0.715 as=0.0798 ps=0.8 w=0.42 l=0.15
X451 a_4993_4175# _023_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X452 VGND a_2957_2999# _088_ VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X453 a_6541_9117# a_6007_8751# a_6446_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.0682 ps=0.745 w=0.42 l=0.15
X454 net10 a_7683_4667# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X455 VGND _013_ a_3677_7497# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X456 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X457 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X459 VGND a_9919_8903# _058_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X460 _089_ a_5177_2487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.33 w=1 l=0.15
X461 a_5411_7815# a_5684_7643# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X462 VPWR _011_ a_4781_9673# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X464 a_7718_6005# a_7550_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.179 ps=1.26 w=0.75 l=0.15
X465 VGND a_5595_8426# _006_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X466 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X467 a_7277_6037# a_7111_6037# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X468 VGND a_8263_6740# _003_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X469 VGND a_2743_7351# net6 VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X470 a_7124_9839# a_6725_9839# a_6998_10205# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X471 _002_ a_6099_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X472 a_4053_6005# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X473 VPWR a_3847_6727# counter\[3\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X474 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X475 a_1475_5461# a_1643_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X476 _061_ a_3243_11293# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.101 ps=0.99 w=0.65 l=0.15
X477 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X478 VGND a_7423_10205# a_7591_10107# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X479 a_5915_5487# counter\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X480 VPWR a_8022_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X481 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X482 VGND a_9983_11195# a_9941_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X483 a_4434_6549# a_4227_6549# a_4610_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0766 ps=0.785 w=0.42 l=0.15
X484 _053_ a_7469_10703# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X485 VGND a_8022_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X486 net3 a_3775_9527# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X487 VPWR _091_ a_2051_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X488 VGND a_5722_6575# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X489 ones[3] a_10239_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X490 VPWR _056_ a_9919_8903# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X492 net10 a_7683_4667# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X493 VGND a_7166_9951# a_7124_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0696 ps=0.765 w=0.42 l=0.15
X494 a_9218_5487# _050_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X495 a_4014_2883# net1 a_3932_2883# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X496 VPWR _032_ a_1499_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X497 a_4864_3829# net6 a_4993_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X498 a_2014_2741# a_1846_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.179 ps=1.26 w=0.75 l=0.15
X499 a_8871_5321# a_8735_5161# a_8451_5175# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
X500 a_4610_6941# a_4363_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X501 VGND a_1407_7119# net2 VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X502 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X503 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X504 _066_ a_9306_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X505 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X506 VGND a_8827_8425# a_8834_8329# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X507 a_3479_7485# a_3259_7497# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.08 w=0.42 l=0.15
X508 _081_ a_6178_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X509 VPWR a_4767_5652# _013_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X510 VGND clknet_1_1__leaf_clk a_6007_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X511 a_8451_5175# a_8735_5161# a_8670_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X512 a_4958_2741# a_4790_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.179 ps=1.26 w=0.75 l=0.15
X513 a_2795_4649# a_2603_4405# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.157 ps=1.17 w=0.42 l=0.15
X514 clknet_1_1__leaf_clk a_8022_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X515 VGND a_9815_11293# a_9983_11195# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X516 VPWR a_5722_6575# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X517 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X518 a_6503_3677# a_5805_3311# a_6246_3423# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X519 VPWR counter\[6\] _078_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X520 a_9815_11293# a_8951_10927# a_9558_11039# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.07 w=0.42 l=0.15
X521 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X522 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X523 a_8022_7119# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X524 clknet_0_clk a_5722_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X525 a_9485_11293# a_8951_10927# a_9390_11293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.0682 ps=0.745 w=0.42 l=0.15
X526 a_8229_9655# _028_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0535 pd=0.675 as=0.122 ps=1.08 w=0.42 l=0.15
X527 VPWR a_2271_2767# a_2439_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X528 VPWR net3 a_9711_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X529 a_7185_2773# a_7019_2773# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X530 a_3081_7119# a_2743_7351# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X531 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X532 a_8447_8439# a_8543_8439# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X533 VGND net7 a_2736_5059# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X534 counter\[6\] a_5751_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X536 counter\[1\] a_1475_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X537 _028_ net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X538 VGND _032_ a_1499_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X539 VGND _037_ a_2695_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X540 _029_ a_3061_9411# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X541 a_9655_9813# net6 a_10136_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.062 ps=0.715 w=0.42 l=0.15
X542 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X543 VGND clknet_1_1__leaf_clk a_7111_6037# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X544 a_6738_9661# a_6423_9527# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X545 VGND net1 _092_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X546 _019_ a_6375_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X547 _048_ a_4627_8320# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.33 w=1 l=0.15
X548 a_5336_2229# _060_ a_5264_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.0535 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X549 VGND a_4053_6005# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X550 a_4363_6575# a_4234_6849# a_3943_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X551 a_3943_6549# a_4234_6849# a_4185_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X552 VPWR a_5215_2767# a_5383_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X553 a_9279_8725# _042_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.312 ps=1.68 w=0.42 l=0.15
X554 _035_ a_6546_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X555 a_3640_6031# _084_ a_3179_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.412 ps=1.82 w=1 l=0.15
X556 VPWR a_9558_11039# a_9485_11293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0766 ps=0.785 w=0.42 l=0.15
X557 VPWR counter\[0\] a_2601_11177# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X559 VGND a_7883_2767# a_8051_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X560 a_3329_6575# counter\[9\] a_3247_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X561 VGND net5 a_9963_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X562 clknet_0_clk a_5722_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X563 a_6997_8751# a_6007_8751# a_6871_9117# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X564 VGND _093_ _011_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X565 VPWR net4 _052_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X566 a_2271_2767# a_1407_2773# a_2014_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.07 w=0.42 l=0.15
X567 VGND a_5722_6575# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X568 a_5722_6575# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X570 a_9919_8903# _055_ a_10153_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X571 VGND a_2014_2741# a_1972_3145# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0696 ps=0.765 w=0.42 l=0.15
X572 _090_ counter\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X573 a_5163_3311# net12 a_4969_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X574 VGND _086_ a_2957_2999# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X575 VGND clknet_0_clk a_8022_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X576 VPWR _008_ a_7357_9673# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X577 a_6527_6263# net11 a_6701_6369# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X578 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X579 VGND _021_ a_9289_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X580 VPWR a_5607_11079# _087_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X581 _024_ net5 a_9043_3561# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X582 a_1846_2767# a_1407_2773# a_1761_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X584 VPWR a_10011_5175# _032_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X585 VGND _000_ a_8369_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X586 VGND _033_ a_5316_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.106 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X587 VGND _054_ a_1867_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X588 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X589 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X590 a_6803_9513# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X591 a_2957_2999# _086_ a_3120_2883# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X592 clknet_1_1__leaf_clk a_8022_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X593 VGND a_5779_5175# _040_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X594 a_1862_5487# a_1475_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X595 VPWR counter\[5\] a_5915_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X596 a_1972_3145# a_1573_2773# a_1846_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X597 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X598 a_2133_6825# net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X599 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X600 VGND a_5411_7815# _076_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X601 VPWR a_4958_2741# a_4885_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0766 ps=0.785 w=0.42 l=0.15
X602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X603 a_7689_4221# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X604 counter\[1\] a_1475_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X605 VPWR clknet_0_clk a_4053_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X606 VGND a_9655_9813# _026_ VGND sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.26 as=0.107 ps=0.98 w=0.65 l=0.15
X607 a_6913_9839# _018_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X608 VGND _033_ a_8352_9527# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X609 a_4227_5161# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X610 _030_ a_2736_5059# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.33 w=1 l=0.15
X611 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X612 clknet_1_1__leaf_clk a_8022_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X613 a_4227_9513# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X614 a_6078_3677# a_5639_3311# a_5993_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X615 VPWR a_4319_7637# a_4326_7937# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X616 VGND _009_ a_4781_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X617 a_3307_9991# _055_ a_3481_9867# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X618 a_2601_11177# counter\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X619 a_9091_5309# a_8871_5321# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.08 w=0.42 l=0.15
X620 a_4885_2767# a_4351_2773# a_4790_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.0682 ps=0.745 w=0.42 l=0.15
X621 a_9827_7351# a_10100_7351# a_10058_7479# VGND sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X622 a_5326_7093# a_5158_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.179 ps=1.26 w=0.75 l=0.15
X623 a_5077_2269# _087_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X624 a_9885_3087# net3 a_10075_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X625 a_6587_3677# a_5805_3311# a_6503_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X627 a_8171_5487# a_7951_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.08 w=0.42 l=0.15
X628 a_5316_5487# net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.106 ps=0.975 w=0.65 l=0.15
X629 a_4909_10089# _092_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X630 VGND _039_ _017_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X631 VPWR a_3307_9991# _080_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X632 a_7111_10383# net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X633 a_7193_10703# _043_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X634 VPWR _042_ a_3801_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X635 a_6204_3311# a_5805_3311# a_6078_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X636 VPWR net7 a_9275_6263# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X637 VGND a_7527_4087# _086_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X638 a_9475_8751# _042_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196 ps=1.33 w=0.42 l=0.15
X639 VPWR counter\[1\] a_1665_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.141 pd=1.32 as=0.0662 ps=0.735 w=0.42 l=0.15
X640 a_6460_5487# _034_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X641 VGND a_4767_5652# _013_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X642 clknet_1_0__leaf_clk a_4053_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X643 a_7515_4765# a_6817_4399# a_7258_4511# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X644 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X645 a_9677_8751# _026_ a_9571_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X646 VGND a_5383_2741# net14 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X647 a_1761_8207# _012_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X648 a_2603_9839# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X649 VPWR a_8022_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X650 a_8022_5461# a_7822_5761# a_8171_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X652 a_9827_7351# a_10100_7351# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X653 _000_ a_8215_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X654 a_3373_6031# _087_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X655 VGND a_8022_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X656 VGND a_7255_3285# _054_ VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X657 a_8815_9527# _044_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.142 ps=1.33 w=0.42 l=0.15
X658 a_2473_6549# net13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.257 ps=1.44 w=0.65 l=0.15
X659 a_9034_8484# a_8834_8329# a_9183_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X660 a_7258_4511# a_7090_4765# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.179 ps=1.26 w=0.75 l=0.15
X661 _020_ a_7847_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X662 VPWR net3 a_10239_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X663 VGND net12 a_3970_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X664 _059_ _058_ a_6013_2473# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X665 _005_ a_6375_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X666 VGND a_6246_3423# a_6204_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0696 ps=0.765 w=0.42 l=0.15
X667 VPWR _068_ _071_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X668 VPWR _074_ a_6009_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X669 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X670 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X671 VPWR _028_ a_8815_9527# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X672 a_4583_5309# a_4363_5321# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.08 w=0.42 l=0.15
X673 a_5126_5487# _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X674 a_1669_6727# _080_ a_1832_6825# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X675 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X676 VPWR a_10075_10357# a_9991_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X677 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X678 VPWR _003_ a_4781_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X679 a_8665_6397# counter\[5\] a_8583_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X680 VGND a_2472_10901# _069_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.172 ps=1.83 w=0.65 l=0.15
X681 a_9728_6147# net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X682 clknet_1_0__leaf_clk a_4053_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X683 VPWR _043_ _046_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X684 VPWR _037_ a_9279_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X685 VPWR a_7423_10205# a_7591_10107# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X686 a_9381_8585# a_8827_8425# a_9034_8484# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X687 _077_ a_9544_3561# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.33 w=1 l=0.15
X688 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X689 counter\[6\] a_5751_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X690 a_3247_6575# counter\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X691 a_5583_7119# a_4719_7125# a_5326_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.07 w=0.42 l=0.15
X692 a_7005_4399# _017_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X693 VGND a_8735_5161# a_8742_5065# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X694 _018_ a_2327_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X695 VPWR a_5722_6575# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X696 VPWR a_2439_8181# net5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X697 VGND a_4227_9513# a_4234_9417# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X698 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X699 a_1941_10749# counter\[2\] a_1841_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X700 a_4418_10927# counter\[3\] a_4322_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X701 a_4351_9839# _049_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X702 VGND a_7815_5461# a_7822_5761# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X703 clknet_0_clk a_5722_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X704 a_8624_10499# counter\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X705 VPWR clk a_5722_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X706 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X707 VPWR _050_ a_4351_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X708 a_5299_2767# a_4517_2773# a_5215_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X709 VGND _059_ a_1748_5303# VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0535 ps=0.675 w=0.42 l=0.15
X710 _000_ a_8215_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X711 a_3148_9655# a_2961_9295# a_3061_9411# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X712 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X713 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X714 VPWR a_8143_6005# a_8059_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X715 a_8785_8207# a_8447_8439# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X716 _075_ a_4338_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X717 a_7515_4765# a_6651_4399# a_7258_4511# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.07 w=0.42 l=0.15
X718 a_8022_5461# a_7815_5461# a_8198_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0766 ps=0.785 w=0.42 l=0.15
X719 VPWR a_9827_7351# _082_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X720 a_5805_3311# a_5639_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X721 a_4864_3829# net5 a_5087_4175# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X722 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X724 VGND clknet_1_0__leaf_clk a_5639_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X725 VPWR _062_ a_9919_8439# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X726 a_9306_7663# counter\[1\] a_9220_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X727 VGND counter\[4\] a_1632_3971# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X728 a_2601_11177# counter\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X729 a_9411_2767# _025_ _012_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X730 VPWR a_5751_7093# a_5667_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X731 VPWR _048_ a_6375_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X732 a_5722_6575# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X734 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X735 a_6013_5309# _034_ a_5941_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X736 VPWR a_4434_6549# a_4363_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.07 w=0.75 l=0.15
X737 VGND a_7039_9019# net7 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X738 _072_ a_1632_3971# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.33 w=1 l=0.15
X739 _051_ a_4351_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X740 VPWR a_1489_4943# a_1589_5059# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X741 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X743 VPWR a_4434_5220# a_4363_5321# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.07 w=0.75 l=0.15
X744 a_4053_6005# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X745 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X746 VPWR _035_ a_8079_9527# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X747 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X748 a_8963_8585# a_8827_8425# a_8543_8439# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
X749 a_5607_11079# counter\[9\] a_5781_10955# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X750 VPWR a_7683_4667# a_7599_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X751 a_7194_5220# a_6987_5161# a_7370_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0766 ps=0.785 w=0.42 l=0.15
X752 _025_ a_9728_6147# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X753 VGND counter\[10\] a_4341_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X754 a_4517_2773# a_4351_2773# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X755 clknet_1_1__leaf_clk a_8022_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X756 a_3215_4551# net8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X757 VGND a_2134_5461# a_2063_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0989 ps=0.995 w=0.64 l=0.15
X758 a_6527_6263# net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X759 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X760 VGND a_9983_11195# net12 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X761 VGND _068_ a_6069_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X762 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X763 a_3330_7396# a_3123_7337# a_3506_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0766 ps=0.785 w=0.42 l=0.15
X764 a_7166_9951# a_6998_10205# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.08 w=0.64 l=0.15
X765 a_7370_4943# a_7123_5321# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X767 VGND a_5215_2767# a_5383_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X768 VPWR a_4053_6005# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X769 VGND a_8143_6005# a_8101_6409# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X770 VGND _084_ a_6989_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X771 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X772 a_3215_4551# net9 a_3389_4427# VGND sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X774 VPWR _060_ a_6835_3968# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X775 a_3506_7119# a_3259_7497# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X776 VPWR a_8355_5175# net4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X777 a_2776_6575# net12 a_2473_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
X778 VPWR a_9279_8725# _043_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X779 a_4719_3311# net11 a_4969_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0877 ps=0.92 w=0.65 l=0.15
X780 a_2014_8181# a_1846_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.179 ps=1.26 w=0.75 l=0.15
X781 clknet_1_1__leaf_clk a_8022_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X782 clknet_0_clk a_5722_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X783 a_4277_8029# a_3939_7815# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X784 VPWR net9 a_10239_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X785 VGND clknet_1_0__leaf_clk a_1407_8213# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X786 VPWR a_7039_9019# net7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X787 VPWR _043_ a_9088_9527# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X788 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X789 VPWR net12 a_9963_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X790 VGND net3 a_10239_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X791 a_10011_5175# _028_ a_10245_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X792 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X793 VPWR clknet_0_clk a_8022_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X794 ready a_8307_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X795 clknet_0_clk a_5722_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X796 VPWR a_3215_4551# _037_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X797 VGND a_4053_6005# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X798 a_9427_9295# net14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X799 a_6725_9839# a_6559_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X800 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X801 a_9551_5652# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X802 a_2695_6144# _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X803 _067_ a_2695_6144# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.33 w=1 l=0.15
X804 VPWR a_1669_6727# _083_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X805 a_10081_8573# _063_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X806 VPWR a_8022_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X807 VPWR _034_ a_5779_5175# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X808 VPWR rst a_1407_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.32 as=0.265 ps=2.53 w=1 l=0.15
X809 a_8583_6397# counter\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X810 clknet_1_0__leaf_clk a_4053_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X811 a_6703_5175# a_6994_5065# a_6945_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X812 VPWR net13 a_7111_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X813 VPWR a_2271_8207# a_2439_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X814 _018_ a_2327_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X815 a_7194_5220# a_6994_5065# a_7343_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X816 a_1714_3971# _068_ a_1632_3971# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X817 VGND a_3775_9527# net3 VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X818 a_3677_7497# a_3130_7241# a_3330_7396# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0682 ps=0.745 w=0.42 l=0.15
X819 a_8762_8573# a_8447_8439# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X820 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X821 ones[4] a_10239_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X822 a_4455_7663# a_4319_7637# a_4035_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
X823 a_6607_5175# a_6703_5175# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X824 a_1927_5461# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X825 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X826 VGND a_2439_8181# net5 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X827 VPWR counter\[1\] _062_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X828 VGND clknet_1_1__leaf_clk a_6651_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X829 a_1841_10749# counter\[3\] a_1769_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X830 ready a_8307_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X831 _002_ a_6099_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X832 _092_ net3 a_2134_4175# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X833 clknet_1_0__leaf_clk a_4053_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X834 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X835 a_7541_5321# a_6987_5161# a_7194_5220# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X836 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X837 a_2271_8207# a_1407_8213# a_2014_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.07 w=0.42 l=0.15
X838 a_9482_10383# a_9043_10389# a_9397_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X839 a_6987_5161# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X840 net12 a_9983_11195# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X842 VGND _090_ a_3368_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X843 VGND a_4043_10901# _068_ VGND sky130_fd_pr__nfet_01v8 ad=0.175 pd=1.26 as=0.107 ps=0.98 w=0.65 l=0.15
X844 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X845 ones[3] a_10239_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X846 a_1761_2767# _007_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X847 a_4338_8751# counter\[4\] a_4252_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X848 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X849 _012_ _024_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.0877 ps=0.92 w=0.65 l=0.15
X850 a_9899_11293# a_9117_10927# a_9815_11293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X851 VGND a_2439_2741# a_2397_3145# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X852 a_5163_3311# net13 _050_ VGND sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.0877 ps=0.92 w=0.65 l=0.15
X853 _044_ a_2736_9001# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.33 w=1 l=0.15
X854 VPWR clknet_0_clk a_4053_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X855 a_6939_9673# a_6803_9513# a_6519_9527# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
X856 a_4781_8573# _046_ a_4709_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X857 a_3970_9839# net12 a_3801_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X858 a_5177_2487# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X859 a_8079_9527# _028_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.142 ps=1.33 w=0.42 l=0.15
X860 a_1573_2773# a_1407_2773# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X861 a_3061_9411# _027_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X862 net8 a_8051_2741# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X863 _091_ net14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X864 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X865 VPWR a_4526_7637# a_4455_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.07 w=0.75 l=0.15
X866 a_7255_3285# a_7431_3285# a_7383_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X867 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X868 a_5595_8426# _079_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X869 VGND _060_ a_3333_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X870 a_9711_2767# _024_ a_9411_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=1.52 w=1 l=0.15
X871 a_9305_10927# _019_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X872 a_3123_7337# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X873 VPWR a_8022_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X874 a_3179_6031# counter\[10\] a_3373_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.412 pd=1.82 as=0.105 ps=1.21 w=1 l=0.15
X875 a_4433_9839# _028_ a_4351_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X876 a_6629_3311# a_5639_3311# a_6503_3677# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X877 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X878 a_4043_10901# counter\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.28 ps=1.62 w=0.42 l=0.15
X879 a_6423_9527# a_6519_9527# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X880 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X881 a_1669_6727# counter\[8\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1 ps=0.985 w=0.42 l=0.15
X882 VPWR _000_ a_8369_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X883 VPWR a_2473_6549# _049_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X884 a_10030_9839# net3 a_9934_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X885 _084_ _080_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X886 a_4969_3311# net11 a_4719_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X887 a_10033_10761# a_9043_10389# a_9907_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X888 VGND net8 a_6546_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X889 a_2839_7351# a_3123_7337# a_3058_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X891 a_2695_4221# _026_ a_2589_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X892 a_2063_5487# a_1927_5461# a_1643_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
X893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X894 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X895 a_6922_5309# a_6607_5175# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X896 VGND net1 a_10075_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X897 VGND _043_ a_2776_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X898 VPWR a_6871_9117# a_7039_9019# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X899 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X900 a_9941_10927# a_8951_10927# a_9815_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X901 VPWR a_4053_6005# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X902 VGND net9 a_10239_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X903 a_8022_7119# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X904 VGND net12 a_9963_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X905 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X906 a_9427_9295# net2 _028_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X907 a_7423_10205# a_6559_9839# a_7166_9951# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.07 w=0.42 l=0.15
X908 VPWR _028_ a_4351_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X909 _024_ net3 a_9126_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X910 a_7093_10205# a_6559_9839# a_6998_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.0682 ps=0.745 w=0.42 l=0.15
X911 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X912 a_9551_5652# _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X913 VPWR _074_ a_5684_7643# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X915 VPWR _010_ a_7541_5321# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X916 _046_ net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X917 VPWR _059_ a_6375_2775# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.32 as=0.166 ps=1.8 w=0.64 l=0.15
X918 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X919 a_2014_2741# a_1846_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.08 w=0.64 l=0.15
X920 VPWR a_9034_8484# a_8963_8585# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.07 w=0.75 l=0.15
X921 VPWR counter\[6\] a_8583_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X922 VPWR a_4053_6005# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X923 _034_ a_2603_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X924 VGND a_6375_2775# _060_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.0877 ps=0.92 w=0.65 l=0.15
X925 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X926 a_9885_3087# net5 _012_ VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0975 ps=0.95 w=0.65 l=0.15
X927 VPWR a_7166_9951# a_7093_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0766 ps=0.785 w=0.42 l=0.15
X928 a_2695_10927# counter\[0\] a_2601_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X929 _074_ a_5915_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X930 _089_ a_5177_2487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X931 VGND a_6671_3579# a_6629_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X932 VPWR _013_ a_3677_7497# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X933 VPWR a_4434_9572# a_4363_9673# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.07 w=0.75 l=0.15
X934 a_2603_4405# _037_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.109 ps=1.36 w=0.42 l=0.15
X935 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X936 a_7465_6031# _002_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X937 a_5997_5487# counter\[5\] a_5915_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X938 VPWR _036_ a_2971_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X939 VPWR _080_ a_10100_7351# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X940 VPWR net7 a_2818_5059# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.33 as=0.0441 ps=0.63 w=0.42 l=0.15
X941 clknet_0_clk a_5722_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X942 a_7626_2741# a_7458_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.179 ps=1.26 w=0.75 l=0.15
X943 ones[4] a_10239_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X944 VPWR a_8022_5461# a_7951_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.07 w=0.75 l=0.15
X945 VPWR _068_ a_5915_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X946 VGND net14 a_3932_2883# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X947 a_9509_6397# net7 a_9437_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X948 VGND a_1547_10004# _007_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X949 VPWR counter\[2\] _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X950 a_5561_7669# _075_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0535 pd=0.675 as=0.122 ps=1.08 w=0.42 l=0.15
X951 a_6917_4221# _060_ a_6835_3968# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X952 VPWR a_8022_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X953 _026_ a_9655_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X954 VGND a_5607_11079# _087_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X955 _050_ _039_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X956 _060_ a_6375_2775# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.32 w=1 l=0.15
X957 _023_ a_3932_2883# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.33 w=1 l=0.15
X958 a_1846_2767# a_1573_2773# a_1761_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X959 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X960 _055_ a_8583_6397# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X961 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X962 VPWR a_1407_7119# net2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X963 VGND net2 a_7431_3285# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X964 a_4885_7125# a_4719_7125# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X965 a_4790_2767# a_4517_2773# a_4705_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X966 a_4043_10901# counter\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0745 pd=0.775 as=0.0777 ps=0.79 w=0.42 l=0.15
X967 a_7005_4399# _017_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X968 a_9397_10383# _020_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X969 a_9390_11293# a_8951_10927# a_9305_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X970 VGND _026_ a_7009_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X971 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X972 a_4162_9661# a_3775_9527# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X973 a_3277_6351# counter\[10\] a_3368_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X974 VGND a_5326_7093# a_5284_7497# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0696 ps=0.765 w=0.42 l=0.15
X975 VGND a_3123_7337# a_3130_7241# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X976 a_6178_9839# counter\[6\] a_6092_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X977 VPWR a_5722_6575# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X978 a_5341_3145# a_4351_2773# a_5215_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X979 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X980 _014_ a_1499_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X981 a_9934_9839# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.175 ps=1.26 w=0.42 l=0.15
X982 a_6614_8863# a_6446_9117# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.08 w=0.64 l=0.15
X983 VGND _076_ a_6375_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X984 _021_ _052_ a_9218_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0959 ps=0.945 w=0.65 l=0.15
X985 VPWR _060_ a_3179_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X986 _063_ a_8624_10499# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X987 a_7883_2767# a_7019_2773# a_7626_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.07 w=0.42 l=0.15
X988 _020_ a_7847_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X989 a_9220_7663# counter\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X990 a_2601_10927# counter\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112 ps=0.995 w=0.65 l=0.15
X991 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X992 VPWR a_4864_3829# _027_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.265 ps=2.53 w=1 l=0.15
X993 a_1643_5461# a_1934_5761# a_1885_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X994 VGND counter\[1\] a_8624_10499# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X995 a_7895_8916# _085_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X996 a_6173_8751# a_6007_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X997 VGND a_7626_2741# a_7584_3145# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0696 ps=0.765 w=0.42 l=0.15
X998 a_4767_5652# _029_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X999 a_2743_7351# a_2839_7351# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1000 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1002 VPWR net11 a_10239_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1003 a_3847_6727# a_3943_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1004 a_4338_8751# counter\[5\] a_4169_9001# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X1005 VGND a_8079_9527# _036_ VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X1006 VPWR clknet_1_1__leaf_clk a_6559_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1007 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1008 clknet_0_clk a_5722_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1009 a_1941_2767# a_1407_2773# a_1846_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.0682 ps=0.745 w=0.42 l=0.15
X1010 _038_ a_2795_4649# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1011 VPWR counter\[8\] _084_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1012 VGND net4 _052_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1013 a_10153_8573# _062_ a_10081_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1015 a_4993_3855# _023_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.172 ps=1.35 w=1 l=0.15
X1016 a_2271_2767# a_1573_2773# a_2014_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1017 VPWR a_2957_2999# _088_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X1018 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1019 a_2961_9295# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1020 a_9046_9655# _028_ a_8965_9655# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0535 ps=0.675 w=0.42 l=0.15
X1021 VGND a_8355_5175# net4 VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1022 clknet_1_0__leaf_clk a_4053_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1023 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1024 _039_ a_2419_4221# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1025 _014_ a_1499_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1026 a_5073_7119# _006_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1027 a_7469_10703# _025_ a_7111_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1028 _050_ net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X1029 VGND a_6527_6263# _042_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1030 a_6078_3677# a_5805_3311# a_5993_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1031 VPWR clknet_0_clk a_8022_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1032 VGND clknet_1_0__leaf_clk a_4719_7125# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1033 VPWR counter\[0\] a_1499_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1034 VGND net5 _024_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1035 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1036 VPWR counter\[4\] a_1714_3971# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.33 as=0.0441 ps=0.63 w=0.42 l=0.15
X1037 VPWR a_7975_6031# a_8143_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1038 a_8827_8425# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1039 VGND a_6503_3677# a_6671_3579# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1040 VGND _031_ a_2795_4649# VGND sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1041 a_7531_5461# a_7815_5461# a_7750_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1042 a_4185_4943# a_3847_5175# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1043 a_2019_2473# _091_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X1044 a_7895_8916# _085_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1045 a_7373_2767# _015_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1046 VPWR _028_ a_5126_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X1047 VGND a_7683_4667# a_7641_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1048 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1049 VGND _051_ a_7847_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1050 a_8543_8439# a_8827_8425# a_8762_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1051 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1053 a_6178_9839# counter\[7\] a_6009_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.138 ps=1.27 w=1 l=0.15
X1054 a_5087_4175# net3 a_4993_4175# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1055 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1056 a_4903_4399# _077_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1057 _053_ a_7469_10703# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.161 ps=1.14 w=0.65 l=0.15
X1058 VPWR a_5583_7119# a_5751_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1059 a_6871_9117# a_6007_8751# a_6614_8863# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.07 w=0.42 l=0.15
X1060 VGND _036_ a_2971_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1061 VPWR a_5722_6575# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1062 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1063 VPWR a_9275_6263# _033_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1064 VGND a_4526_7637# a_4455_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0989 ps=0.995 w=0.64 l=0.15
X1065 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1066 a_7277_6037# a_7111_6037# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1067 _079_ a_4903_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.33 w=1 l=0.15
X1068 a_9655_9813# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0745 pd=0.775 as=0.0777 ps=0.79 w=0.42 l=0.15
X1069 VGND a_3847_5175# counter\[9\] VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1070 net14 a_5383_2741# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1071 a_6614_8863# a_6446_9117# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.179 ps=1.26 w=0.75 l=0.15
X1072 VPWR a_6246_3423# a_6173_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0766 ps=0.785 w=0.42 l=0.15
X1073 a_6607_5175# a_6703_5175# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1074 a_3847_6727# a_3943_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1075 VGND _047_ a_4781_8573# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1076 a_9390_11293# a_9117_10927# a_9305_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1077 a_7383_3311# _058_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.101 ps=0.99 w=0.42 l=0.15
X1078 net8 a_8051_2741# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1079 a_6725_9839# a_6559_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1080 a_2051_6575# _040_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1081 clknet_1_1__leaf_clk a_8022_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1082 VPWR a_9650_10357# a_9577_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0766 ps=0.785 w=0.42 l=0.15
X1083 VPWR _028_ a_3061_9411# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.0744 ps=0.815 w=0.42 l=0.15
X1084 a_4363_5321# a_4227_5161# a_3943_5175# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
X1085 a_2355_2767# a_1573_2773# a_2271_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1086 VPWR a_9815_11293# a_9983_11195# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1087 a_6173_3677# a_5639_3311# a_6078_3677# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.0682 ps=0.745 w=0.42 l=0.15
X1088 VPWR net5 a_9711_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X1089 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1090 a_7009_5487# net7 _031_ VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1091 VGND a_3307_9991# _080_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1093 a_5057_4399# _077_ a_4985_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1094 a_4035_7637# a_4319_7637# a_4254_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1095 a_3943_5175# a_4227_5161# a_4162_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1096 VPWR a_7718_6005# a_7645_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0766 ps=0.785 w=0.42 l=0.15
X1097 a_2472_10901# counter\[1\] a_2695_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X1098 _092_ net1 a_2051_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1099 a_8310_9655# _035_ a_8229_9655# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0535 ps=0.675 w=0.42 l=0.15
X1100 VPWR net1 a_2019_2473# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.35 as=0.16 ps=1.32 w=1 l=0.15
X1101 a_6377_5737# _023_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1102 VGND _088_ a_5336_2229# VGND sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.08 as=0.0535 ps=0.675 w=0.42 l=0.15
X1103 VPWR net6 a_2603_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1104 VPWR net6 a_10239_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1105 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1106 clknet_1_0__leaf_clk a_4053_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1107 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1108 a_5642_7669# _060_ a_5561_7669# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0535 ps=0.675 w=0.42 l=0.15
X1109 a_1761_8207# _012_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1110 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1111 a_7645_6031# a_7111_6037# a_7550_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.0682 ps=0.745 w=0.42 l=0.15
X1112 VPWR a_8022_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1113 net13 a_10075_10357# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1114 a_7111_10383# net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1115 net1 a_1407_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.162 ps=1.32 w=1 l=0.15
X1116 a_2014_8181# a_1846_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.08 w=0.64 l=0.15
X1117 VGND a_8022_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1118 VGND _058_ _059_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1119 a_9815_11293# a_9117_10927# a_9558_11039# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1120 a_7773_5853# a_7363_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1121 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1122 VPWR _084_ a_6835_3968# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X1123 VPWR clknet_1_0__leaf_clk a_4351_2773# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1124 _093_ a_1925_2473# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.172 ps=1.35 w=1 l=0.15
X1125 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1126 a_6987_5161# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1127 VGND _053_ _021_ VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1128 a_2375_10615# _060_ a_2609_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1129 a_3330_7396# a_3130_7241# a_3479_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1130 a_4252_8751# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1131 a_1573_8213# a_1407_8213# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1132 VGND _066_ a_2849_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1133 VPWR net12 _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.135 ps=1.27 w=1 l=0.15
X1134 a_4767_5652# _029_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1135 a_4053_6005# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1136 a_2481_5487# a_1934_5761# a_2134_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0682 ps=0.745 w=0.42 l=0.15
X1137 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1138 VPWR counter\[0\] a_3063_11293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.109 ps=1.36 w=0.42 l=0.15
X1139 a_7090_4765# a_6651_4399# a_7005_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1140 VGND a_1475_5461# counter\[1\] VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X1141 _077_ a_9544_3561# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1142 a_5077_2269# _087_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1143 VPWR _060_ a_5411_7815# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0744 ps=0.815 w=0.42 l=0.15
X1144 VGND net11 a_10239_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1145 VPWR counter\[10\] a_3247_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X1146 VGND a_2014_8181# a_1972_8585# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0696 ps=0.765 w=0.42 l=0.15
X1147 a_4627_8320# _046_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1148 _056_ a_1665_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.141 ps=1.32 w=1 l=0.15
X1149 VGND a_5722_6575# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1150 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1151 a_1573_2773# a_1407_2773# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1152 a_8079_5162# _073_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1153 _016_ a_5126_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1154 a_3677_7497# a_3123_7337# a_3330_7396# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1155 a_4319_7637# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1156 ones[0] a_10239_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1157 VGND a_4319_7637# a_4326_7937# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1158 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1159 VPWR a_5722_6575# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1160 VPWR a_5779_5175# _040_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1161 a_1846_8207# a_1407_8213# a_1761_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1162 a_10011_5175# _028_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1163 VGND a_7039_9019# a_6997_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1164 a_7216_4399# a_6817_4399# a_7090_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1165 a_8451_5175# a_8742_5065# a_8693_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1166 VPWR a_4053_6005# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1167 _085_ a_6835_3968# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1168 a_6945_4943# a_6607_5175# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1170 a_7951_5487# a_7815_5461# a_7531_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
X1171 VGND a_2271_2767# a_2439_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1172 VGND net14 _091_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1173 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1174 a_1769_10749# a_1499_10383# a_1665_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1176 a_9608_10761# a_9209_10389# a_9482_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1177 _057_ a_3247_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.33 w=1 l=0.15
X1178 VPWR a_7431_3285# a_7255_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1179 a_1972_8585# a_1573_8213# a_1846_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1181 _047_ a_3970_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X1182 VGND a_7258_4511# a_7216_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0696 ps=0.765 w=0.42 l=0.15
X1183 VPWR _090_ a_3640_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X1184 _078_ _074_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1185 a_9977_7479# _081_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0535 pd=0.675 as=0.122 ps=1.08 w=0.42 l=0.15
X1186 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1187 a_2375_10615# _072_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.33 w=0.42 l=0.15
X1188 VPWR net14 a_8307_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1189 VGND a_7975_6031# a_8143_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1190 a_6803_9513# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1191 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1192 a_6989_4221# _083_ a_6917_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1193 a_7431_3285# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X1194 a_2419_4221# _026_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1195 a_4043_10901# counter\[1\] a_4524_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.062 ps=0.715 w=0.42 l=0.15
X1196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1197 VGND a_8447_8439# counter\[5\] VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1198 a_8059_6031# a_7277_6037# a_7975_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1199 a_5997_6351# counter\[1\] _065_ VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1201 VGND a_8942_5220# a_8871_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0989 ps=0.995 w=0.64 l=0.15
X1202 a_7815_5461# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1203 a_2736_5059# _026_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1204 clknet_1_0__leaf_clk a_4053_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1205 a_7619_8916# _089_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1206 VGND net11 a_2736_9001# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1207 VPWR a_9983_11195# a_9899_11293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1208 a_3801_10089# _040_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1209 a_3401_6575# counter\[8\] a_3329_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1210 a_6519_9527# a_6803_9513# a_6738_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1211 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1212 VPWR a_7527_4087# _086_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1213 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1214 VGND a_9907_10383# a_10075_10357# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1215 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1216 VPWR net3 a_2603_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1217 VGND a_5583_7119# a_5751_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1218 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1219 a_7289_10703# net12 a_7193_10703# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.107 ps=0.98 w=0.65 l=0.15
X1220 a_9626_3561# _074_ a_9544_3561# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1221 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1223 a_5667_7119# a_4885_7125# a_5583_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1224 a_2019_2473# net2 a_1925_2473# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X1225 a_4227_9513# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1226 _011_ _092_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1228 a_9919_8903# _057_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.33 w=0.42 l=0.15
X1229 VGND _011_ a_4781_9673# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1231 a_4969_3311# net12 a_5163_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1232 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1233 VGND a_4958_2741# a_4916_3145# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0696 ps=0.765 w=0.42 l=0.15
X1234 a_3943_9527# a_4227_9513# a_4162_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1235 a_6761_9295# a_6423_9527# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1236 VPWR counter\[4\] a_8583_6397# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1238 _052_ net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1239 a_2501_4221# net10 a_2419_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1240 VGND _025_ _012_ VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1241 VGND net14 a_8307_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1242 a_2839_7351# a_3130_7241# a_3081_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1243 a_7507_10205# a_6725_9839# a_7423_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1244 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1245 a_7363_5461# a_7531_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1246 _041_ _040_ a_2133_6825# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1247 VGND a_7194_5220# a_7123_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0989 ps=0.995 w=0.64 l=0.15
X1248 VPWR a_3847_5175# counter\[9\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1249 VPWR net10 a_10239_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1250 VPWR a_7039_9019# a_6955_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1251 a_7599_4765# a_6817_4399# a_7515_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1252 VGND _048_ a_6375_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1253 VGND _068_ a_6089_9615# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1254 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1255 _051_ a_4351_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.33 w=1 l=0.15
X1256 VGND net6 a_10239_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1257 a_2593_2473# _041_ _017_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1258 a_1846_8207# a_1573_8213# a_1761_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1259 a_7619_8916# _089_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1260 VPWR a_4053_6005# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1261 a_10136_9839# net5 a_10030_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.062 pd=0.715 as=0.0798 ps=0.8 w=0.42 l=0.15
X1262 clknet_0_clk a_5722_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1263 a_5805_3311# a_5639_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1264 VPWR a_5722_6575# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1265 VPWR a_6803_9513# a_6810_9417# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1266 a_3259_7497# a_3130_7241# a_2839_7351# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1267 clknet_1_1__leaf_clk a_8022_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1268 a_9118_4943# a_8871_5321# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1269 a_2743_7351# a_2839_7351# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1270 a_7761_4221# _055_ a_7689_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1271 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1272 a_2603_9839# net7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1273 VPWR _050_ a_9135_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X1274 a_1861_6351# counter\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1275 VGND counter\[2\] a_9306_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X1276 a_4185_9295# a_3775_9527# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1277 a_9397_10383# _020_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1278 VPWR _066_ a_2695_6144# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X1279 a_8263_6740# _070_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1280 VGND clknet_0_clk a_4053_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1281 a_1589_5059# _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X1282 a_4583_9661# a_4363_9673# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.08 w=0.42 l=0.15
X1283 a_8079_5162# _073_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1284 VGND a_5751_7093# a_5709_7497# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1285 VGND a_6871_9117# a_7039_9019# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1286 a_8079_9527# a_8352_9527# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.108 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1287 a_4705_2767# _022_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1289 a_4993_3855# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1290 VPWR clknet_1_1__leaf_clk a_9043_10389# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1291 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1292 clknet_1_0__leaf_clk a_4053_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1293 ones[5] a_10239_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1294 VPWR net14 a_4014_2883# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.33 as=0.0441 ps=0.63 w=0.42 l=0.15
X1295 VGND _010_ a_7541_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1296 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1297 ones[0] a_10239_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1298 a_6092_9839# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1299 clknet_0_clk a_5722_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1300 a_3939_7815# a_4035_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1301 VPWR net11 a_6527_6263# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X1302 VGND clk a_5722_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1303 a_8871_5321# a_8742_5065# a_8451_5175# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1304 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1305 a_2773_9839# net6 a_2685_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1306 a_9289_5321# a_8742_5065# a_8942_5220# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0682 ps=0.745 w=0.42 l=0.15
X1307 a_2472_10901# counter\[3\] a_2601_11177# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1308 VGND net3 a_2879_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1309 a_1941_8207# a_1407_8213# a_1846_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.0682 ps=0.745 w=0.42 l=0.15
X1310 a_4363_9673# a_4227_9513# a_3943_9527# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
X1311 clknet_1_0__leaf_clk a_4053_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1312 a_7527_4087# counter\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1313 a_7363_5461# a_7531_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1314 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1315 net14 a_5383_2741# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X1316 VPWR a_9919_8903# _058_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1317 ones[10] a_8307_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1318 a_10081_8751# _057_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X1319 VGND counter\[0\] a_1499_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1320 VPWR clknet_1_1__leaf_clk a_7019_2773# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1321 VPWR a_5722_6575# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1322 VPWR _037_ a_2419_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1323 _071_ counter\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1324 a_9516_10927# a_9117_10927# a_9390_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1325 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1326 VGND _008_ a_7357_9673# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1327 a_6817_4399# a_6651_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1328 a_9289_5321# a_8735_5161# a_8942_5220# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1329 a_7343_5309# a_7123_5321# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.08 w=0.42 l=0.15
X1330 a_6246_3423# a_6078_3677# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.179 ps=1.26 w=0.75 l=0.15
X1331 a_1489_4943# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1332 a_6246_3423# a_6078_3677# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.08 w=0.64 l=0.15
X1333 VPWR a_9983_11195# net12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1334 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1335 VGND a_6423_9527# counter\[8\] VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1336 a_7123_5321# a_6994_5065# a_6703_5175# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1337 clknet_1_1__leaf_clk a_8022_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1338 _070_ a_1589_5059# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122 ps=1.08 w=0.65 l=0.15
X1339 a_4781_5321# a_4234_5065# a_4434_5220# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0682 ps=0.745 w=0.42 l=0.15
X1340 VPWR counter\[9\] a_3247_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1341 a_8079_9527# a_8352_9527# a_8310_9655# VGND sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1343 ones[1] a_9963_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1344 a_8735_5161# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1345 a_5434_5737# _033_ a_5126_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.162 pd=1.32 as=0.22 ps=1.44 w=1 l=0.15
X1346 a_8101_6409# a_7111_6037# a_7975_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1347 VPWR _061_ a_8215_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1348 a_3939_7815# a_4035_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1349 VGND a_4434_6549# a_4363_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0989 ps=0.995 w=0.64 l=0.15
X1350 a_8706_10499# counter\[0\] a_8624_10499# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1351 VPWR _076_ a_6375_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1352 counter\[0\] a_7363_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1353 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1354 VGND _043_ a_9088_9527# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.108 ps=1.36 w=0.42 l=0.15
X1355 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1356 VGND _025_ a_7469_10703# VGND sky130_fd_pr__nfet_01v8 ad=0.161 pd=1.14 as=0.184 ps=1.21 w=0.65 l=0.15
X1357 VPWR a_5411_7815# _076_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1358 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1359 a_1665_10383# a_1499_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X1360 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1361 VGND net10 a_10239_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1362 VGND a_2271_8207# a_2439_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1363 _066_ a_9306_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X1364 a_10011_5175# _031_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.33 w=0.42 l=0.15
X1365 VGND net14 _028_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0877 ps=0.92 w=0.65 l=0.15
X1366 a_7159_9661# a_6939_9673# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.08 w=0.42 l=0.15
X1367 a_2355_8207# a_1573_8213# a_2271_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1368 a_9544_3561# _074_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1371 VGND _001_ a_2481_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1372 VGND a_5722_6575# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1373 a_7626_2741# a_7458_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.08 w=0.64 l=0.15
X1374 VPWR a_4227_6549# a_4234_6849# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1375 _010_ a_3179_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.0877 ps=0.92 w=0.65 l=0.15
X1376 VPWR _045_ a_2327_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1377 _078_ counter\[6\] a_9589_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1378 a_9650_10357# a_9482_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.08 w=0.64 l=0.15
X1379 a_3943_6549# a_4227_6549# a_4162_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1380 a_7385_10703# net13 a_7289_10703# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1381 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1382 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1383 a_2818_9001# _039_ a_2736_9001# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1384 a_2397_3145# a_1407_2773# a_2271_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1385 VPWR net9 a_5434_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.162 ps=1.32 w=1 l=0.15
X1386 a_6093_6351# counter\[0\] a_5997_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.107 ps=0.98 w=0.65 l=0.15
X1387 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1388 a_9991_10383# a_9209_10389# a_9907_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1389 a_5595_8426# _079_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1390 VGND _061_ a_8215_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1391 a_9655_9813# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.28 ps=1.62 w=0.42 l=0.15
X1392 _025_ a_9728_6147# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.33 w=1 l=0.15
X1393 a_8263_6740# _070_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1394 a_4053_6005# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1395 VPWR a_7194_5220# a_7123_5321# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.07 w=0.75 l=0.15
X1396 VPWR a_4227_5161# a_4234_5065# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1397 a_2051_3855# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.148 ps=1.29 w=1 l=0.15
X1398 VGND a_9919_8439# _064_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1399 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1400 VPWR _034_ a_6377_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1401 _035_ a_6546_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.257 ps=1.44 w=0.65 l=0.15
X1402 a_8543_8439# a_8834_8329# a_8785_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1403 ones[5] a_10239_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1404 a_8670_5309# a_8355_5175# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1405 VPWR a_4053_6005# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1406 clknet_0_clk a_5722_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1407 VPWR a_6503_3677# a_6671_3579# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1408 VPWR net3 a_9655_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X1409 VPWR net3 a_2019_2473# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1410 a_9411_2767# _024_ a_9711_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1411 VPWR _059_ a_1589_5059# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.0744 ps=0.815 w=0.42 l=0.15
X1412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1413 VPWR _051_ a_7847_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1414 a_2691_6825# net13 a_2473_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1415 a_7750_5487# a_7363_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1416 clknet_1_1__leaf_clk a_8022_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0578 ps=0.695 w=0.42 l=0.15
X1417 a_9810_6147# net2 a_9728_6147# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1418 a_7641_4399# a_6651_4399# a_7515_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1419 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1420 a_5722_6575# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1421 VPWR counter\[1\] a_8706_10499# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.33 as=0.0441 ps=0.63 w=0.42 l=0.15
X1422 net12 a_9983_11195# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1423 a_5411_7815# _075_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.142 ps=1.33 w=0.42 l=0.15
X1424 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1425 a_4341_4399# counter\[9\] _090_ VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1426 a_2283_5487# a_2063_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.121 ps=1.08 w=0.42 l=0.15
X1427 VGND clknet_1_0__leaf_clk a_4351_2773# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1428 a_4526_7637# a_4319_7637# a_4702_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0766 ps=0.785 w=0.42 l=0.15
X1429 counter\[0\] a_7363_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1430 net11 a_7591_10107# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1431 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1432 VGND a_2439_8181# a_2397_8585# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1433 a_9117_10927# a_8951_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1434 a_2877_4649# a_2603_4405# a_2795_4649# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1435 VGND a_4053_6005# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1436 VGND counter\[10\] a_3401_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1437 a_3333_10927# a_3063_11293# a_3243_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.109 ps=1.36 w=0.42 l=0.15
X1438 VGND _039_ a_4719_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1440 VPWR a_8447_8439# counter\[5\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1441 a_9919_8903# _055_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1442 a_3389_4427# net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.112 ps=1.04 w=0.42 l=0.15
X1443 VGND a_4227_6549# a_4234_6849# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1444 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1445 VPWR a_8815_9527# _045_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1446 a_5607_11079# _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X1447 a_10075_3087# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1448 a_4702_8029# a_4455_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1449 VPWR counter\[6\] a_9626_3561# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.33 as=0.0441 ps=0.63 w=0.42 l=0.15
X1450 a_2134_5461# a_1934_5761# a_2283_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1451 VPWR a_3775_9527# net3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1452 VPWR a_1407_10927# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1453 a_9919_8439# _063_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.33 w=0.42 l=0.15
X1454 VPWR _028_ _041_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X1455 a_7258_4511# a_7090_4765# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.08 w=0.64 l=0.15
X1456 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1457 ones[9] a_8583_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1458 clknet_0_clk a_5722_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1459 a_5326_7093# a_5158_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.121 ps=1.08 w=0.64 l=0.15
X1460 VPWR net14 a_9427_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1461 a_9117_10927# a_8951_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1462 a_1547_10004# _082_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1463 VPWR a_1927_5461# a_1934_5761# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1464 _034_ a_2603_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X1465 VPWR _060_ a_2695_6144# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1466 a_5583_7119# a_4885_7125# a_5326_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1467 a_4185_6941# a_3847_6727# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.111 ps=1.37 w=0.42 l=0.15
X1468 VGND net10 a_2051_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.107 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1469 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1470 VPWR a_7010_9572# a_6939_9673# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.109 ps=1.07 w=0.75 l=0.15
X1471 a_2481_5487# a_1927_5461# a_2134_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1472 clknet_1_0__leaf_clk a_4053_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1473 a_2777_6397# _060_ a_2695_6144# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1474 VGND a_8022_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1475 a_7166_9951# a_6998_10205# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.179 ps=1.26 w=0.75 l=0.15
X1476 a_4254_7663# a_3939_7815# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X1477 VPWR net7 a_9279_8725# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X1478 a_2965_10703# _080_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1479 ones[1] a_9963_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1480 a_6173_8751# a_6007_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1481 a_9711_2767# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1482 _012_ net5 a_9885_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1483 VPWR _039_ a_2593_2473# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1484 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1485 a_3884_9839# _042_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.172 ps=1.83 w=0.65 l=0.15
X1486 a_2609_10749# _071_ a_2537_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1487 a_9907_10383# a_9043_10389# a_9650_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.07 w=0.42 l=0.15
X1488 a_7883_2767# a_7185_2773# a_7626_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1489 a_9137_7913# counter\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X1490 a_9577_10383# a_9043_10389# a_9482_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.0682 ps=0.745 w=0.42 l=0.15
X1491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1492 a_4873_7663# a_4326_7937# a_4526_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0682 ps=0.745 w=0.42 l=0.15
X1493 a_3932_2883# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1494 a_7550_6031# a_7277_6037# a_7465_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1495 counter\[7\] a_2439_2741# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1496 a_7527_4087# counter\[8\] a_7761_4221# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1497 VGND clknet_1_1__leaf_clk a_9043_10389# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1498 a_3307_9991# _068_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.167 ps=1.39 w=0.42 l=0.15
X1499 ones[9] a_8583_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1500 VPWR a_9551_5652# _001_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1501 VPWR a_1475_5461# counter\[1\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1502 VGND net2 _028_ VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X1503 _068_ a_4043_10901# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X1504 a_6013_2473# net2 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1505 VPWR a_2375_10615# _073_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1506 a_7527_4087# _068_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.33 w=0.42 l=0.15
X1507 VPWR a_4053_6005# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1508 clknet_1_1__leaf_clk a_8022_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1509 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1510 a_4363_6575# a_4227_6549# a_3943_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
X1511 VPWR _039_ _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1512 VPWR a_6375_2775# _060_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1513 a_2134_5461# a_1927_5461# a_2310_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0766 ps=0.785 w=0.42 l=0.15
X1514 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1515 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1516 a_5779_5175# _023_ a_6013_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1517 VPWR counter\[10\] _090_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1518 _050_ net13 a_5163_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X1519 VGND _045_ a_2327_9295# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1520 a_9827_7351# _081_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0744 pd=0.815 as=0.142 ps=1.33 w=0.42 l=0.15
X1521 _048_ a_4627_8320# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1522 a_5073_7119# _006_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.109 ps=1.36 w=0.42 l=0.15
X1523 a_1676_5303# a_1489_4943# a_1589_5059# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.108 ps=1.36 w=0.42 l=0.15
X1524 net1 a_1407_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0682 ps=0.745 w=0.42 l=0.15
X1525 VGND clknet_0_clk a_4053_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1526 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1527 a_2375_10615# _060_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1528 VPWR a_6987_5161# a_6994_5065# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1529 ones[7] a_10239_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1530 a_3368_6351# _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1531 VPWR a_5077_2269# a_5177_2487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X1532 a_4505_9839# _049_ a_4433_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1533 a_2310_5853# a_2063_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0766 pd=0.785 as=0.179 ps=1.26 w=0.42 l=0.15
X1534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1535 VPWR clknet_1_0__leaf_clk a_1407_2773# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1536 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1537 a_5316_5487# _038_ a_5216_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.114 ps=1 w=0.65 l=0.15
X1538 VGND a_4434_9572# a_4363_9673# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0989 ps=0.995 w=0.64 l=0.15
X1539 a_6998_10205# a_6559_9839# a_6913_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1540 a_2211_2223# _091_ a_2115_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.107 ps=0.98 w=0.65 l=0.15
X1541 VPWR a_8827_8425# a_8834_8329# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1542 a_10173_5309# _031_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.132 ps=1.14 w=0.42 l=0.15
X1543 a_5779_5175# _037_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.142 ps=1.33 w=0.42 l=0.15
X1544 a_9381_8585# a_8834_8329# a_9034_8484# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0682 ps=0.745 w=0.42 l=0.15
X1545 VPWR a_2961_9295# a_3061_9411# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.108 ps=1.36 w=0.42 l=0.15
X1546 VPWR net12 a_2691_6825# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1547 VGND counter\[7\] a_6178_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.257 pd=1.44 as=0.0894 ps=0.925 w=0.65 l=0.15
X1548 VGND a_5722_6575# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1549 a_2134_4175# _091_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0959 pd=0.945 as=0.172 ps=1.83 w=0.65 l=0.15
X1550 clknet_0_clk a_5722_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.138 ps=1.27 w=1 l=0.15
X1551 _075_ a_4338_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1552 a_10153_8751# _056_ a_10081_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1553 a_7967_2767# a_7185_2773# a_7883_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1554 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1555 VPWR a_6423_9527# counter\[8\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1556 a_4781_9673# a_4234_9417# a_4434_9572# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0578 pd=0.695 as=0.0682 ps=0.745 w=0.42 l=0.15
X1557 VPWR a_7515_4765# a_7683_4667# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1558 VGND clk a_5722_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1559 VGND net6 a_4864_3829# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.107 ps=0.98 w=0.65 l=0.15
X1560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1561 a_5158_7119# a_4719_7125# a_5073_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1562 VGND a_9279_8725# _043_ VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X1563 VPWR a_2014_2741# a_1941_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.179 pd=1.26 as=0.0766 ps=0.785 w=0.42 l=0.15
X1564 VPWR clknet_1_1__leaf_clk a_7111_6037# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X1565 VGND a_7718_6005# a_7676_6409# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0696 ps=0.765 w=0.42 l=0.15
X1566 VPWR _060_ a_3243_11293# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.228 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1567 a_2063_5487# a_1934_5761# a_1643_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1568 VPWR _023_ a_9043_3561# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.29 as=0.265 ps=2.53 w=1 l=0.15
X1569 a_6939_9673# a_6810_9417# a_6519_9527# VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1570 a_9279_8725# net7 a_9677_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X1571 VGND a_4053_6005# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1573 a_7458_2767# a_7019_2773# a_7373_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1574 VPWR a_5595_8426# _006_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1575 a_7423_10205# a_6725_9839# a_7166_9951# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1576 a_5284_7497# a_4885_7125# a_5158_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1577 VGND a_8022_5461# a_7951_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.121 pd=1.08 as=0.0989 ps=0.995 w=0.64 l=0.15
X1578 _028_ net2 a_9427_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1579 VGND a_7515_4765# a_7683_4667# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1580 _029_ a_3061_9411# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.33 w=1 l=0.15
X1581 VGND net1 a_2211_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X1582 a_10075_3087# net3 a_9885_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.0877 pd=0.92 as=0.0877 ps=0.92 w=0.65 l=0.15
X1583 a_5722_6575# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
X1584 a_4885_7125# a_4719_7125# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1585 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1586 counter\[2\] a_8143_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1587 net2 a_1407_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0682 ps=0.745 w=0.42 l=0.15
X1588 VPWR a_7591_10107# a_7507_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1589 a_10058_7479# _060_ a_9977_7479# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0535 ps=0.675 w=0.42 l=0.15
X1590 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1591 net9 a_6671_3579# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1592 a_8753_6397# counter\[4\] a_8665_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1594 a_7584_3145# a_7185_2773# a_7458_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1595 VGND counter\[6\] a_8859_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1596 VGND a_4053_6005# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1597 a_9275_6263# net8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1598 VGND _067_ a_6099_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1599 VPWR a_9907_10383# a_10075_10357# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1600 VPWR a_8051_2741# a_7967_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.111 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1601 VPWR _060_ a_4903_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1602 a_9209_10389# a_9043_10389# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1603 VPWR _071_ a_2375_10615# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X1604 _093_ a_1925_2473# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.172 pd=1.83 as=0.112 ps=0.995 w=0.65 l=0.15
X1605 VPWR a_8022_7119# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1606 VGND _005_ a_9381_8585# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1607 a_3970_9839# _040_ a_3884_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1608 a_9275_6263# net8 a_9509_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1609 a_7465_6031# _002_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1610 _039_ a_2419_4221# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X1611 _084_ counter\[8\] a_2965_10703# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0877 ps=0.92 w=0.65 l=0.15
X1612 a_6955_9117# a_6173_8751# a_6871_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1613 VPWR _004_ a_4873_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0578 ps=0.695 w=0.42 l=0.15
X1614 VGND net7 a_10239_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1616 a_6913_9839# _018_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.109 ps=1.36 w=0.42 l=0.15
X1617 VGND clknet_1_1__leaf_clk a_7019_2773# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1618 a_2271_8207# a_1573_8213# a_2014_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1619 a_2961_9295# _026_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.108 pd=1.36 as=0.109 ps=1.36 w=0.42 l=0.15
X1620 ones[2] a_10239_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1621 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1622 VPWR _047_ a_4627_8320# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.33 as=0.0662 ps=0.735 w=0.42 l=0.15
X1623 VGND a_9551_5652# _001_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1624 VPWR net7 a_2419_4221# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1625 a_8583_6397# counter\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1626 a_6703_5175# a_6987_5161# a_6922_5309# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1627 _044_ a_2736_9001# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1628 VGND a_10011_5175# _032_ VGND sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1629 clknet_1_0__leaf_clk a_4053_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1630 VGND a_8022_7119# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1631 VGND net14 a_9728_6147# VGND sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1632 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1633 VPWR net3 a_4993_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1634 a_6009_10089# counter\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.138 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
D2 VGND net6 sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06 area=4.347e+11
X1635 a_5158_7119# a_4885_7125# a_5073_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0682 pd=0.745 as=0.0578 ps=0.695 w=0.42 l=0.15
X1636 a_7975_6031# a_7277_6037# a_7718_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1637 a_8735_5161# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1638 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1639 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1640 _019_ a_6375_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1641 a_7815_5461# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1642 clknet_0_clk a_5722_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1643 VGND a_3215_4551# _037_ VGND sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1644 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1645 ones[7] a_10239_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
C0 net11 net3 0.421f
C1 net13 net6 1.43f
C2 _014_ _039_ 0.173f
C3 _093_ _054_ 0.436f
C4 _002_ a_7277_6037# 0.195f
C5 _052_ counter\[7\] 2.18f
C6 _088_ net2 0.671f
C7 _062_ _074_ 0.339f
C8 _010_ a_6994_5065# 0.569f
C9 _045_ _033_ 0.114f
C10 VPWR a_4338_8751# 0.204f
C11 a_5326_7093# a_4719_7125# 0.141f
C12 _062_ counter\[9\] 0.383f
C13 _004_ counter\[0\] 0.517f
C14 VPWR a_3243_11293# 0.169f
C15 a_6651_4399# a_7258_4511# 0.138f
C16 net1 a_2439_2741# 0.115f
C17 a_6810_9417# clknet_1_1__leaf_clk 0.207f
C18 net8 counter\[10\] 0.34f
C19 a_8942_5220# VPWR 0.244f
C20 counter\[7\] _034_ 0.574f
C21 _004_ counter\[8\] 0.149f
C22 a_5722_6575# counter\[2\] 0.268f
C23 counter\[1\] a_8624_10499# 0.199f
C24 net8 _023_ 0.186f
C25 _078_ net7 0.358f
C26 _043_ _033_ 0.124f
C27 _039_ _017_ 0.11f
C28 _074_ counter\[0\] 0.267f
C29 net7 net3 0.249f
C30 _093_ _011_ 0.12f
C31 net6 _039_ 0.118f
C32 a_7531_5461# VPWR 0.184f
C33 net13 _086_ 0.376f
C34 _028_ a_4351_9839# 0.213f
C35 VPWR a_4363_6575# 0.174f
C36 _058_ net2 1.07f
C37 _019_ net14 0.132f
C38 _003_ a_8263_6740# 0.109f
C39 a_6939_9673# a_6803_9513# 0.141f
C40 a_8834_8329# a_8963_8585# 0.117f
C41 _014_ _087_ 0.151f
C42 net8 _025_ 1.48f
C43 a_4434_9572# a_4363_9673# 0.24f
C44 net5 _092_ 0.19f
C45 _001_ VPWR 1.02f
C46 _032_ counter\[4\] 0.743f
C47 counter\[6\] _037_ 1.5f
C48 _043_ _082_ 0.499f
C49 _068_ _044_ 0.325f
C50 VPWR _047_ 0.276f
C51 _084_ _040_ 0.268f
C52 VPWR a_7626_2741# 0.174f
C53 ones[1] a_9963_2223# 0.111f
C54 a_2375_10615# _072_ 0.198f
C55 counter\[9\] counter\[8\] 0.328f
C56 _022_ a_1867_9295# 0.109f
C57 _028_ a_9088_9527# 0.126f
C58 _031_ _034_ 0.252f
C59 _037_ clknet_1_1__leaf_clk 0.963f
C60 a_4363_5321# VPWR 0.178f
C61 VPWR a_2014_8181# 0.222f
C62 net9 a_10239_6575# 0.194f
C63 a_6913_9839# _018_ 0.113f
C64 VPWR a_9650_10357# 0.174f
C65 a_1407_8213# a_1846_8207# 0.273f
C66 _064_ VPWR 0.417f
C67 net4 net11 0.719f
C68 _087_ _017_ 0.344f
C69 net11 _042_ 0.151f
C70 VPWR a_2971_3311# 0.264f
C71 VPWR a_3943_6549# 0.178f
C72 _067_ a_6099_4399# 0.193f
C73 a_6651_4399# VPWR 0.446f
C74 a_3215_4551# net8 0.162f
C75 a_9728_6147# net14 0.175f
C76 a_7277_6037# counter\[4\] 0.453f
C77 _053_ counter\[0\] 0.709f
C78 _026_ _037_ 0.506f
C79 counter\[1\] clknet_0_clk 0.585f
C80 net13 net1 0.461f
C81 _025_ _028_ 0.664f
C82 _048_ _076_ 0.121f
C83 ones[4] _028_ 0.166f
C84 _085_ clknet_1_1__leaf_clk 0.299f
C85 VPWR a_5684_7643# 0.161f
C86 _005_ _085_ 0.303f
C87 net6 _015_ 0.138f
C88 a_2971_3311# _036_ 0.206f
C89 _028_ _060_ 0.123f
C90 a_3847_5175# counter\[9\] 0.113f
C91 _071_ counter\[4\] 0.115f
C92 VPWR a_2271_2767# 0.216f
C93 _045_ _044_ 0.105f
C94 net8 _002_ 0.2f
C95 net4 net7 0.441f
C96 net7 _042_ 0.347f
C97 counter\[1\] a_1665_10383# 0.181f
C98 VPWR a_4767_5652# 0.207f
C99 _068_ _043_ 0.603f
C100 _086_ _087_ 0.24f
C101 net14 _023_ 0.15f
C102 a_5383_2741# a_5215_2767# 0.311f
C103 VPWR a_7847_10383# 0.206f
C104 a_1665_10383# counter\[3\] 0.165f
C105 net1 _039_ 0.595f
C106 _053_ _050_ 0.142f
C107 net14 _025_ 0.248f
C108 net11 a_6725_9839# 0.212f
C109 VPWR counter\[5\] 1.37f
C110 _043_ _044_ 0.317f
C111 VPWR counter\[6\] 1.83f
C112 counter\[2\] _037_ 0.243f
C113 VPWR a_3259_7497# 0.2f
C114 _084_ _055_ 0.12f
C115 net14 _060_ 0.141f
C116 a_6671_3579# a_6503_3677# 0.311f
C117 a_6614_8863# a_6173_8751# 0.111f
C118 _077_ _060_ 0.112f
C119 _009_ _042_ 0.551f
C120 ones[8] ones[9] 0.122f
C121 VPWR clknet_1_1__leaf_clk 5.12f
C122 counter\[9\] _068_ 0.449f
C123 a_6559_9839# clknet_1_1__leaf_clk 0.259f
C124 _005_ VPWR 0.603f
C125 a_8827_8425# clknet_1_1__leaf_clk 0.466f
C126 net5 _027_ 0.159f
C127 a_4319_7637# VPWR 0.479f
C128 _069_ counter\[2\] 0.357f
C129 _005_ a_8827_8425# 0.133f
C130 VPWR a_5751_7093# 0.395f
C131 counter\[5\] net10 0.38f
C132 VPWR a_1643_5461# 0.201f
C133 clknet_1_0__leaf_clk a_5639_3311# 0.219f
C134 counter\[6\] net10 0.269f
C135 _086_ a_2957_2999# 0.1f
C136 a_6607_5175# a_6703_5175# 0.311f
C137 _021_ _074_ 0.325f
C138 VPWR _026_ 2.56f
C139 _055_ ones[9] 0.109f
C140 _072_ net3 0.178f
C141 VPWR a_5583_7119# 0.184f
C142 VPWR a_3932_2883# 0.18f
C143 VPWR clknet_1_0__leaf_clk 5.65f
C144 clknet_0_clk a_5722_6575# 1.69f
C145 _001_ _050_ 0.38f
C146 _066_ _028_ 1.02f
C147 a_9827_7351# _060_ 0.101f
C148 ones[5] VPWR 0.31f
C149 VPWR a_9907_10383# 0.174f
C150 net9 net4 0.93f
C151 a_3247_6575# counter\[10\] 0.196f
C152 _066_ _035_ 0.146f
C153 VPWR _076_ 0.44f
C154 _012_ clknet_1_0__leaf_clk 0.24f
C155 _008_ a_7357_9673# 0.115f
C156 _010_ _004_ 0.159f
C157 VPWR counter\[7\] 1.76f
C158 _077_ _002_ 0.189f
C159 _028_ _040_ 0.192f
C160 _026_ a_2961_9295# 0.142f
C161 a_2795_4649# a_2603_4405# 0.101f
C162 VPWR a_10011_5175# 0.234f
C163 _062_ counter\[6\] 0.142f
C164 clknet_1_0__leaf_clk _036_ 0.317f
C165 a_2375_10615# _060_ 0.17f
C166 _026_ net10 0.405f
C167 VPWR a_5126_5487# 0.419f
C168 a_2736_9001# _039_ 0.102f
C169 clknet_1_0__leaf_clk net10 0.118f
C170 _032_ _092_ 0.69f
C171 net7 net2 0.467f
C172 a_5411_7815# a_5684_7643# 0.168f
C173 _066_ net14 0.166f
C174 _026_ _059_ 0.11f
C175 _053_ _021_ 0.176f
C176 a_8735_5161# a_8942_5220# 0.26f
C177 a_3123_7337# VPWR 0.709f
C178 _058_ _085_ 0.368f
C179 a_4719_7125# clknet_1_0__leaf_clk 0.25f
C180 VPWR counter\[2\] 2.63f
C181 _002_ a_6375_4399# 0.121f
C182 VPWR _031_ 2.37f
C183 _070_ counter\[2\] 0.219f
C184 VPWR a_9558_11039# 0.176f
C185 _070_ _031_ 0.113f
C186 _004_ _074_ 0.431f
C187 counter\[9\] _043_ 0.259f
C188 _076_ _059_ 0.116f
C189 counter\[1\] _020_ 0.193f
C190 _016_ _040_ 0.142f
C191 _028_ counter\[4\] 0.232f
C192 a_6939_9673# a_7010_9572# 0.24f
C193 _008_ a_6810_9417# 0.262f
C194 net12 net5 0.173f
C195 net8 _055_ 1.24f
C196 _001_ _068_ 0.357f
C197 _041_ _039_ 0.846f
C198 VPWR _088_ 1.36f
C199 counter\[0\] clknet_1_1__leaf_clk 0.302f
C200 counter\[5\] _033_ 1.3f
C201 VPWR a_9275_6263# 0.203f
C202 _026_ _080_ 0.289f
C203 net11 _034_ 0.643f
C204 a_4326_7937# a_4455_7663# 0.119f
C205 counter\[8\] clknet_1_1__leaf_clk 0.16f
C206 a_9983_11195# a_9815_11293# 0.311f
C207 _065_ clknet_1_0__leaf_clk 0.473f
C208 _049_ _028_ 0.883f
C209 a_1925_2473# net1 0.124f
C210 a_6607_5175# VPWR 0.398f
C211 VPWR a_2439_8181# 0.453f
C212 _014_ a_6173_8751# 0.181f
C213 _050_ counter\[5\] 0.113f
C214 VPWR a_7255_3285# 0.157f
C215 a_7019_2773# a_7626_2741# 0.136f
C216 clknet_1_1__leaf_clk _033_ 0.236f
C217 _057_ a_9919_8903# 0.215f
C218 _053_ _043_ 0.316f
C219 counter\[1\] _056_ 0.138f
C220 _080_ counter\[7\] 0.476f
C221 _027_ _087_ 0.191f
C222 VPWR a_4227_6549# 0.441f
C223 _031_ _059_ 0.151f
C224 net8 net6 0.152f
C225 _001_ _021_ 0.148f
C226 _026_ counter\[8\] 0.992f
C227 _073_ a_8079_5162# 0.188f
C228 _039_ a_2419_4221# 0.111f
C229 VPWR _058_ 1.91f
C230 net13 net12 1.22f
C231 clknet_1_0__leaf_clk counter\[8\] 0.296f
C232 _082_ clknet_1_1__leaf_clk 0.787f
C233 clknet_0_clk _037_ 0.641f
C234 a_4781_9673# a_4234_9417# 0.102f
C235 _050_ clknet_1_1__leaf_clk 0.403f
C236 a_4234_5065# net12 0.247f
C237 net7 _034_ 0.114f
C238 clk _003_ 0.182f
C239 _012_ _058_ 0.105f
C240 _026_ _033_ 0.163f
C241 _078_ counter\[10\] 0.142f
C242 _062_ counter\[2\] 0.329f
C243 counter\[6\] _024_ 0.117f
C244 net9 net2 0.126f
C245 _093_ _040_ 0.347f
C246 counter\[10\] net3 0.399f
C247 VPWR a_4227_9513# 0.439f
C248 _081_ _018_ 0.231f
C249 a_6810_9417# net11 0.121f
C250 net5 _022_ 0.238f
C251 net1 ones[9] 0.162f
C252 _019_ net4 0.171f
C253 _023_ net3 0.767f
C254 counter\[8\] counter\[7\] 0.124f
C255 _073_ VPWR 1.06f
C256 _073_ _070_ 0.236f
C257 a_8143_6005# a_7975_6031# 0.311f
C258 _054_ net2 2.01f
C259 _026_ _050_ 1.2f
C260 _025_ net3 0.369f
C261 clknet_1_0__leaf_clk _050_ 0.263f
C262 counter\[7\] _033_ 0.165f
C263 a_10239_2223# net3 0.201f
C264 VPWR a_8624_10499# 0.148f
C265 _078_ _060_ 0.876f
C266 counter\[2\] counter\[0\] 1.57f
C267 _072_ counter\[3\] 0.448f
C268 _060_ net3 0.379f
C269 counter\[2\] a_9306_7663# 0.186f
C270 a_5126_5487# _033_ 0.111f
C271 net14 _055_ 0.183f
C272 _068_ counter\[5\] 1.09f
C273 _001_ a_9551_5652# 0.135f
C274 a_3943_5175# a_4234_5065# 0.192f
C275 a_6246_3423# a_5639_3311# 0.136f
C276 net11 _037_ 0.217f
C277 _050_ counter\[7\] 0.381f
C278 net12 a_9117_10927# 0.12f
C279 VPWR a_5607_11079# 0.233f
C280 net13 _022_ 0.143f
C281 _062_ a_4227_6549# 0.464f
C282 counter\[7\] a_6178_9839# 0.178f
C283 VPWR a_7718_6005# 0.194f
C284 a_2019_2473# VPWR 0.211f
C285 VPWR a_6246_3423# 0.185f
C286 _062_ _058_ 0.582f
C287 a_8735_5161# clknet_1_1__leaf_clk 0.316f
C288 _053_ _063_ 0.82f
C289 VPWR ones[10] 0.273f
C290 a_3063_11293# _060_ 0.124f
C291 _005_ _068_ 0.34f
C292 VPWR a_1407_2773# 0.771f
C293 net14 net6 0.593f
C294 _048_ net7 0.282f
C295 _064_ a_9551_5652# 0.183f
C296 VPWR a_1927_5461# 0.727f
C297 VPWR _008_ 0.461f
C298 net9 _034_ 0.23f
C299 counter\[2\] _089_ 0.496f
C300 net7 _037_ 0.41f
C301 clknet_1_1__leaf_clk a_7019_2773# 0.256f
C302 VPWR a_6099_4399# 0.258f
C303 _091_ clknet_1_0__leaf_clk 0.146f
C304 _068_ _026_ 0.569f
C305 VPWR clknet_0_clk 3.06f
C306 VPWR a_4517_2773# 0.282f
C307 net4 _023_ 0.451f
C308 _073_ _080_ 0.143f
C309 _021_ clknet_1_1__leaf_clk 0.104f
C310 net4 _025_ 0.557f
C311 _066_ ones[6] 0.105f
C312 ones[4] net4 0.203f
C313 net1 a_1407_10927# 0.173f
C314 _079_ clknet_1_0__leaf_clk 1.38f
C315 a_9381_8585# _005_ 0.115f
C316 net14 _086_ 0.826f
C317 rst net2 0.103f
C318 net4 _060_ 0.146f
C319 VPWR a_1665_10383# 0.367f
C320 _016_ _086_ 0.642f
C321 _019_ a_9305_10927# 0.115f
C322 _026_ a_9655_9813# 0.114f
C323 clknet_0_clk net10 0.249f
C324 _074_ a_5684_7643# 0.123f
C325 _092_ _028_ 0.292f
C326 _045_ clknet_1_1__leaf_clk 0.456f
C327 VPWR a_2473_6549# 0.21f
C328 a_4363_5321# a_4227_5161# 0.136f
C329 counter\[0\] a_8624_10499# 0.117f
C330 _022_ _087_ 0.111f
C331 _040_ net3 0.4f
C332 a_3061_9411# _028_ 0.217f
C333 _093_ _017_ 0.107f
C334 net12 _038_ 0.245f
C335 a_2601_11177# VPWR 0.201f
C336 net6 _093_ 0.202f
C337 a_8742_5065# a_8871_5321# 0.119f
C338 a_3330_7396# VPWR 0.267f
C339 a_9650_10357# a_9482_10383# 0.24f
C340 VPWR net11 1.85f
C341 net6 a_2603_9839# 0.159f
C342 _068_ counter\[2\] 1.15f
C343 _067_ counter\[10\] 0.509f
C344 VPWR a_4790_2767# 0.245f
C345 VPWR a_8215_8751# 0.208f
C346 _060_ a_6375_2775# 0.158f
C347 _043_ clknet_1_1__leaf_clk 0.245f
C348 _073_ _082_ 0.232f
C349 _074_ counter\[5\] 0.239f
C350 _062_ clknet_0_clk 0.975f
C351 _073_ _050_ 0.211f
C352 a_7822_5761# _000_ 0.195f
C353 _073_ _089_ 0.237f
C354 _074_ counter\[6\] 2.09f
C355 _004_ clknet_1_1__leaf_clk 0.316f
C356 _013_ net12 0.438f
C357 counter\[1\] _025_ 0.551f
C358 _010_ clknet_1_0__leaf_clk 0.153f
C359 a_9728_6147# net2 0.123f
C360 net1 net14 0.349f
C361 ones[4] ones[3] 0.111f
C362 a_4526_7637# a_4455_7663# 0.24f
C363 a_4319_7637# _004_ 0.139f
C364 clknet_0_clk _080_ 0.13f
C365 net11 net10 0.294f
C366 _067_ _060_ 0.104f
C367 _084_ net12 0.538f
C368 VPWR ones[1] 0.142f
C369 _026_ _043_ 0.113f
C370 VPWR net7 5.76f
C371 counter\[1\] _060_ 0.554f
C372 _070_ net7 0.111f
C373 clknet_1_0__leaf_clk _043_ 0.165f
C374 a_8022_7119# _081_ 0.135f
C375 VPWR a_9544_3561# 0.15f
C376 a_8447_8439# a_8543_8439# 0.311f
C377 clknet_0_clk counter\[0\] 0.188f
C378 counter\[3\] _060_ 0.146f
C379 net13 net5 0.148f
C380 _066_ net4 0.243f
C381 _049_ net3 0.1f
C382 _053_ a_7847_10383# 0.116f
C383 a_2603_4405# _037_ 0.17f
C384 net9 _085_ 0.657f
C385 _026_ _074_ 0.194f
C386 _023_ net2 0.673f
C387 _025_ a_7469_10703# 0.168f
C388 net7 net10 0.202f
C389 VPWR a_2743_7351# 0.432f
C390 net6 a_10239_3311# 0.221f
C391 _053_ counter\[6\] 0.391f
C392 VPWR a_4434_9572# 0.243f
C393 _025_ net2 0.122f
C394 counter\[9\] _026_ 0.138f
C395 VPWR _009_ 0.546f
C396 _015_ a_7185_2773# 0.279f
C397 VPWR a_10239_5487# 0.252f
C398 clknet_1_0__leaf_clk counter\[9\] 0.5f
C399 _010_ _031_ 0.362f
C400 a_1573_8213# VPWR 0.345f
C401 _018_ _028_ 0.926f
C402 counter\[7\] _074_ 0.292f
C403 a_8834_8329# _028_ 0.172f
C404 net7 _059_ 0.152f
C405 _092_ _093_ 0.231f
C406 _053_ clknet_1_1__leaf_clk 0.75f
C407 _012_ a_1573_8213# 0.281f
C408 _043_ counter\[2\] 0.409f
C409 _055_ net3 0.32f
C410 net1 _093_ 0.104f
C411 _063_ clknet_1_1__leaf_clk 0.131f
C412 a_10239_9295# net11 0.203f
C413 counter\[5\] a_4338_8751# 0.171f
C414 _043_ _031_ 0.175f
C415 _084_ _022_ 0.117f
C416 net11 counter\[0\] 0.132f
C417 _004_ _031_ 0.339f
C418 a_7683_4667# a_7515_4765# 0.311f
C419 _027_ _028_ 0.388f
C420 VPWR _020_ 0.245f
C421 _016_ a_5805_3311# 0.261f
C422 counter\[8\] net11 0.204f
C423 a_4227_5161# clknet_1_0__leaf_clk 0.224f
C424 net13 a_10075_10357# 0.136f
C425 _052_ _023_ 0.11f
C426 VPWR net9 2.33f
C427 counter\[2\] _074_ 0.887f
C428 counter\[1\] _066_ 0.825f
C429 net9 _070_ 0.406f
C430 _080_ net7 0.602f
C431 net11 _033_ 0.16f
C432 _025_ _052_ 0.849f
C433 a_5595_8426# _006_ 0.109f
C434 VPWR a_5177_2487# 0.207f
C435 a_5077_2269# VPWR 0.17f
C436 VPWR a_6671_3579# 0.398f
C437 net6 net3 1.39f
C438 net4 _051_ 0.222f
C439 _001_ counter\[6\] 0.102f
C440 counter\[9\] counter\[2\] 0.19f
C441 counter\[9\] _031_ 0.516f
C442 VPWR _054_ 0.79f
C443 _082_ net11 0.161f
C444 _034_ _023_ 0.246f
C445 _046_ _028_ 1.1f
C446 a_9711_2767# net3 0.103f
C447 net8 net12 0.316f
C448 net9 _036_ 0.442f
C449 a_6725_9839# a_7166_9951# 0.119f
C450 net11 _050_ 0.185f
C451 VPWR a_2014_2741# 0.213f
C452 counter\[8\] net7 1.29f
C453 VPWR _056_ 1.61f
C454 a_5073_7119# _006_ 0.131f
C455 a_2695_6144# VPWR 0.222f
C456 a_8051_2741# a_7883_2767# 0.311f
C457 a_7895_8916# _085_ 0.188f
C458 VPWR _029_ 0.52f
C459 _069_ rst 0.249f
C460 a_7277_6037# a_7111_6037# 0.962f
C461 a_4903_4399# _060_ 0.176f
C462 a_8079_9527# _028_ 0.226f
C463 a_2063_5487# a_1934_5761# 0.127f
C464 a_2134_5461# a_1927_5461# 0.273f
C465 a_4227_5161# _031_ 0.443f
C466 _008_ _044_ 0.159f
C467 VPWR _011_ 0.301f
C468 _086_ net3 0.142f
C469 VPWR pulse 0.238f
C470 _053_ counter\[2\] 0.215f
C471 _001_ _026_ 0.316f
C472 net4 _055_ 0.209f
C473 _042_ _055_ 0.24f
C474 _001_ clknet_1_0__leaf_clk 0.111f
C475 _019_ _085_ 0.107f
C476 _064_ clknet_1_1__leaf_clk 0.109f
C477 counter\[1\] counter\[4\] 0.393f
C478 VPWR a_3307_9991# 0.2f
C479 VPWR _072_ 0.824f
C480 _018_ _093_ 0.101f
C481 a_6651_4399# clknet_1_1__leaf_clk 0.31f
C482 a_6614_8863# a_6007_8751# 0.136f
C483 a_3943_9527# a_4234_9417# 0.192f
C484 counter\[0\] _020_ 0.224f
C485 _068_ net11 0.903f
C486 VPWR a_7895_8916# 0.211f
C487 VPWR a_8143_6005# 0.381f
C488 _092_ net3 0.168f
C489 VPWR a_5215_2767# 0.18f
C490 _009_ _050_ 0.23f
C491 _023_ _037_ 0.47f
C492 net1 net3 0.892f
C493 a_1846_2767# a_1407_2773# 0.273f
C494 rst VPWR 0.262f
C495 _056_ _080_ 0.128f
C496 _079_ net11 0.34f
C497 net14 net12 0.16f
C498 ones[3] a_10239_4399# 0.111f
C499 counter\[1\] _014_ 0.307f
C500 a_2481_5487# a_1934_5761# 0.102f
C501 _019_ VPWR 0.699f
C502 counter\[5\] clknet_1_1__leaf_clk 0.178f
C503 clk _093_ 1.29f
C504 net9 _033_ 0.284f
C505 _084_ net5 0.209f
C506 a_6527_6263# net11 0.134f
C507 counter\[6\] clknet_1_1__leaf_clk 0.308f
C508 _015_ _039_ 0.819f
C509 net8 _000_ 0.123f
C510 _068_ net7 0.706f
C511 _037_ _060_ 0.223f
C512 clknet_0_clk _043_ 0.108f
C513 a_2736_5059# _030_ 0.107f
C514 a_4885_7125# net14 0.466f
C515 _072_ a_1632_3971# 0.123f
C516 net9 _050_ 0.19f
C517 _005_ clknet_1_1__leaf_clk 0.164f
C518 _026_ counter\[5\] 0.227f
C519 a_6614_8863# a_6446_9117# 0.24f
C520 _080_ a_3307_9991# 0.115f
C521 a_7515_4765# a_6817_4399# 0.195f
C522 _063_ a_8624_10499# 0.105f
C523 VPWR a_4351_9839# 0.18f
C524 clknet_0_clk _074_ 0.166f
C525 a_3215_4551# _037_ 0.12f
C526 _003_ a_4234_6849# 0.184f
C527 a_4363_6575# a_4227_6549# 0.136f
C528 VPWR a_9728_6147# 0.159f
C529 _021_ net7 0.17f
C530 a_6803_9513# a_6810_9417# 0.969f
C531 _055_ net2 0.125f
C532 _026_ clknet_1_1__leaf_clk 0.611f
C533 _072_ counter\[0\] 0.131f
C534 _056_ _082_ 0.11f
C535 counter\[7\] counter\[5\] 0.22f
C536 VPWR a_9815_11293# 0.185f
C537 counter\[7\] counter\[6\] 0.349f
C538 VPWR a_9088_9527# 0.167f
C539 a_4319_7637# clknet_1_0__leaf_clk 0.224f
C540 _007_ a_1573_2773# 0.234f
C541 a_5583_7119# a_5751_7093# 0.311f
C542 VPWR a_8447_8439# 0.427f
C543 ones[0] ones[1] 0.16f
C544 _079_ _009_ 1.34f
C545 counter\[7\] clknet_1_1__leaf_clk 0.203f
C546 a_8815_9527# _028_ 0.121f
C547 a_6519_9527# a_6423_9527# 0.311f
C548 VPWR counter\[10\] 0.728f
C549 clknet_1_0__leaf_clk _026_ 0.125f
C550 _064_ _058_ 1.13f
C551 VPWR _023_ 0.907f
C552 net2 _017_ 0.499f
C553 _034_ _051_ 0.822f
C554 ones[2] ones[1] 0.103f
C555 counter\[2\] counter\[5\] 0.37f
C556 _010_ net7 1.36f
C557 a_6503_3677# a_5805_3311# 0.192f
C558 net11 _074_ 0.302f
C559 a_3123_7337# a_3259_7497# 0.141f
C560 _072_ _082_ 0.292f
C561 clknet_1_0__leaf_clk _076_ 1.38f
C562 VPWR a_7683_4667# 0.415f
C563 _066_ _037_ 0.724f
C564 VPWR _025_ 1.29f
C565 rst counter\[0\] 0.306f
C566 _026_ counter\[7\] 0.4f
C567 ones[4] VPWR 0.299f
C568 VPWR a_10239_2223# 0.216f
C569 _043_ net7 0.3f
C570 _019_ counter\[0\] 0.196f
C571 VPWR a_5595_8426# 0.279f
C572 _007_ _093_ 0.154f
C573 clknet_1_0__leaf_clk counter\[7\] 0.783f
C574 _027_ net3 0.44f
C575 counter\[10\] _036_ 0.143f
C576 counter\[2\] clknet_1_1__leaf_clk 0.126f
C577 _012_ _025_ 0.224f
C578 _031_ clknet_1_1__leaf_clk 0.725f
C579 VPWR _060_ 7.02f
C580 VPWR a_2327_9295# 0.212f
C581 _041_ net3 0.106f
C582 a_9043_10389# a_9209_10389# 0.969f
C583 a_7166_9951# a_6998_10205# 0.24f
C584 _013_ _087_ 0.306f
C585 _012_ _060_ 0.205f
C586 _034_ _055_ 0.117f
C587 net7 _074_ 0.159f
C588 _025_ net10 0.29f
C589 a_3123_7337# clknet_1_0__leaf_clk 0.261f
C590 _026_ _031_ 0.303f
C591 _023_ _059_ 0.489f
C592 a_3215_4551# VPWR 0.216f
C593 clk net3 0.175f
C594 _074_ a_9544_3561# 0.109f
C595 counter\[9\] net7 0.363f
C596 net10 _060_ 1.41f
C597 a_3179_6031# _060_ 0.123f
C598 _058_ counter\[6\] 0.695f
C599 net12 a_3970_9839# 0.176f
C600 counter\[2\] counter\[7\] 0.117f
C601 _091_ _072_ 0.276f
C602 a_9275_6263# _026_ 0.206f
C603 _059_ _060_ 0.365f
C604 _057_ _035_ 0.273f
C605 _031_ a_10011_5175# 0.202f
C606 _068_ a_3307_9991# 0.162f
C607 a_7373_2767# a_7185_2773# 0.102f
C608 a_6835_3968# _060_ 0.167f
C609 _058_ clknet_1_1__leaf_clk 0.379f
C610 VPWR _002_ 1.06f
C611 _005_ _058_ 0.165f
C612 a_9983_11195# net12 0.177f
C613 a_6614_8863# VPWR 0.197f
C614 _088_ counter\[7\] 0.19f
C615 _062_ _060_ 0.136f
C616 a_2839_7351# a_3130_7241# 0.195f
C617 _069_ counter\[4\] 0.215f
C618 VPWR a_6803_9513# 0.659f
C619 _050_ a_4351_9839# 0.216f
C620 a_4227_6549# clknet_1_0__leaf_clk 0.217f
C621 _073_ clknet_1_1__leaf_clk 0.118f
C622 VPWR a_8583_6397# 0.417f
C623 VPWR _066_ 1.12f
C624 _056_ _045_ 2.75f
C625 _080_ _060_ 1.65f
C626 net12 net3 0.866f
C627 _057_ net14 0.125f
C628 a_6817_4399# a_7258_4511# 0.116f
C629 _025_ counter\[0\] 0.252f
C630 a_7815_5461# a_8022_5461# 0.273f
C631 _002_ net10 0.225f
C632 a_1846_2767# a_2014_2741# 0.24f
C633 net11 _047_ 0.21f
C634 clknet_1_0__leaf_clk a_4227_9513# 0.671f
C635 VPWR _040_ 0.773f
C636 counter\[0\] _060_ 0.289f
C637 _070_ _040_ 0.238f
C638 _073_ _026_ 0.19f
C639 _056_ _043_ 0.111f
C640 VPWR a_7166_9951# 0.183f
C641 counter\[8\] _060_ 1.03f
C642 a_6725_9839# _018_ 0.227f
C643 a_7166_9951# a_6559_9839# 0.136f
C644 a_7822_5761# net8 0.482f
C645 _066_ net10 0.827f
C646 VPWR a_7883_2767# 0.196f
C647 a_7550_6031# a_7111_6037# 0.26f
C648 _050_ _023_ 0.129f
C649 net13 a_9043_10389# 0.447f
C650 a_3939_7815# counter\[4\] 0.137f
C651 net1 _052_ 0.175f
C652 _007_ net3 0.43f
C653 _025_ _082_ 0.317f
C654 _073_ counter\[7\] 0.495f
C655 ones[10] clknet_1_1__leaf_clk 0.164f
C656 _001_ net7 0.138f
C657 _083_ _072_ 0.928f
C658 _032_ _030_ 0.334f
C659 _040_ net10 0.222f
C660 _039_ _028_ 0.124f
C661 _082_ _060_ 0.293f
C662 net13 net14 0.195f
C663 _055_ _085_ 0.123f
C664 VPWR counter\[4\] 4.39f
C665 _022_ net3 0.84f
C666 _008_ clknet_1_1__leaf_clk 0.178f
C667 _050_ _060_ 0.173f
C668 a_7423_10205# a_6725_9839# 0.192f
C669 _084_ _071_ 0.338f
C670 VPWR a_6817_4399# 0.314f
C671 counter\[1\] a_4053_6005# 0.278f
C672 VPWR _051_ 2.25f
C673 a_7465_6031# _002_ 0.127f
C674 net5 _093_ 0.117f
C675 a_6559_9839# _051_ 0.423f
C676 VPWR _049_ 0.775f
C677 _066_ _080_ 0.624f
C678 clknet_1_0__leaf_clk a_1407_2773# 0.307f
C679 _062_ _040_ 0.3f
C680 VPWR ones[8] 0.242f
C681 clknet_1_0__leaf_clk a_1927_5461# 0.25f
C682 a_8834_8329# a_8543_8439# 0.195f
C683 net10 counter\[4\] 0.308f
C684 _086_ _037_ 0.24f
C685 _058_ a_7255_3285# 0.202f
C686 VPWR a_3801_10089# 0.267f
C687 _080_ _040_ 0.221f
C688 VPWR a_7123_5321# 0.202f
C689 clknet_1_0__leaf_clk a_4517_2773# 0.287f
C690 net11 counter\[5\] 0.21f
C691 _066_ a_9306_7663# 0.119f
C692 _068_ _023_ 0.142f
C693 net11 counter\[6\] 0.765f
C694 _036_ _049_ 0.162f
C695 a_3130_7241# _013_ 0.255f
C696 a_3330_7396# a_3259_7497# 0.24f
C697 _066_ counter\[8\] 0.121f
C698 a_1573_8213# a_2014_8181# 0.119f
C699 VPWR a_10239_4399# 0.254f
C700 net8 _038_ 0.149f
C701 VPWR _014_ 1.42f
C702 VPWR _055_ 3.7f
C703 net11 clknet_1_1__leaf_clk 0.389f
C704 _001_ net9 1.65f
C705 VPWR a_8263_6740# 0.269f
C706 _068_ _060_ 0.306f
C707 a_8263_6740# _070_ 0.205f
C708 _061_ _081_ 0.424f
C709 a_1499_6031# _014_ 0.108f
C710 _086_ _085_ 0.158f
C711 counter\[4\] a_1632_3971# 0.203f
C712 a_7005_4399# _017_ 0.118f
C713 a_1407_8213# VPWR 0.757f
C714 _066_ _082_ 0.142f
C715 counter\[1\] net12 1.7f
C716 _065_ counter\[4\] 0.406f
C717 a_5595_8426# _079_ 0.197f
C718 _026_ net11 0.221f
C719 VPWR _017_ 1.87f
C720 a_1407_8213# _012_ 0.135f
C721 clknet_1_0__leaf_clk net11 0.194f
C722 VPWR net6 4.97f
C723 net8 _084_ 1.18f
C724 counter\[6\] a_9544_3561# 0.17f
C725 clknet_0_clk counter\[2\] 0.139f
C726 net12 counter\[3\] 0.772f
C727 net7 clknet_1_1__leaf_clk 0.341f
C728 ones[6] a_10239_7663# 0.11f
C729 counter\[0\] counter\[4\] 0.76f
C730 _018_ _034_ 0.204f
C731 _028_ _038_ 0.152f
C732 VPWR a_9711_2767# 0.512f
C733 _043_ a_9088_9527# 0.132f
C734 VPWR a_8022_5461# 0.25f
C735 net11 counter\[7\] 0.103f
C736 _010_ counter\[10\] 0.168f
C737 _047_ _029_ 0.213f
C738 _069_ net1 0.106f
C739 ones[0] a_10239_2223# 0.11f
C740 _009_ counter\[5\] 0.24f
C741 _083_ _023_ 0.153f
C742 VPWR a_4864_3829# 0.191f
C743 a_10239_9295# ones[8] 0.125f
C744 _062_ _055_ 0.132f
C745 _026_ net7 1.6f
C746 counter\[4\] _033_ 0.423f
C747 clk a_5722_6575# 0.311f
C748 clknet_1_0__leaf_clk net7 0.294f
C749 VPWR _086_ 3.39f
C750 _043_ _023_ 0.19f
C751 counter\[8\] _049_ 0.221f
C752 a_7039_9019# VPWR 0.488f
C753 _070_ _086_ 0.169f
C754 _045_ a_2327_9295# 0.199f
C755 a_9919_8439# VPWR 0.22f
C756 _014_ _080_ 0.148f
C757 _080_ _055_ 0.12f
C758 _009_ clknet_1_1__leaf_clk 0.191f
C759 a_3123_7337# a_3330_7396# 0.273f
C760 _059_ _017_ 0.297f
C761 a_7847_10383# _020_ 0.114f
C762 VPWR a_7010_9572# 0.271f
C763 net6 _059_ 0.136f
C764 _012_ _086_ 0.113f
C765 counter\[2\] net11 0.273f
C766 _025_ _043_ 0.325f
C767 _083_ _060_ 0.347f
C768 _050_ counter\[4\] 0.902f
C769 net5 net3 3.86f
C770 a_7373_2767# _015_ 0.115f
C771 a_7258_4511# a_7090_4765# 0.24f
C772 _014_ counter\[0\] 0.14f
C773 a_7123_5321# a_6994_5065# 0.111f
C774 a_8022_5461# a_7951_5487# 0.24f
C775 _086_ _036_ 0.16f
C776 a_9963_9295# VPWR 0.196f
C777 net9 counter\[5\] 0.121f
C778 net9 counter\[6\] 0.21f
C779 _014_ counter\[8\] 0.104f
C780 counter\[10\] counter\[9\] 0.239f
C781 a_9827_7351# _081_ 0.202f
C782 _050_ _049_ 0.186f
C783 ones[8] _082_ 0.151f
C784 _068_ _040_ 1.32f
C785 _004_ _060_ 0.594f
C786 _025_ _074_ 0.253f
C787 net5 a_9963_2223# 0.205f
C788 a_1573_8213# clknet_1_0__leaf_clk 0.235f
C789 _020_ clknet_1_1__leaf_clk 0.208f
C790 a_8951_10927# a_9117_10927# 0.964f
C791 VPWR a_7591_10107# 0.388f
C792 _055_ _033_ 0.362f
C793 net9 clknet_1_1__leaf_clk 0.108f
C794 VPWR a_6987_5161# 0.464f
C795 VPWR _092_ 1.92f
C796 a_4767_5652# _029_ 0.198f
C797 _031_ net7 0.555f
C798 a_8583_10927# ready 0.109f
C799 VPWR net1 6.47f
C800 VPWR a_3061_9411# 0.2f
C801 net13 net3 0.213f
C802 _012_ _092_ 1.81f
C803 _082_ _055_ 1.67f
C804 _054_ clknet_1_1__leaf_clk 0.277f
C805 a_7039_9019# a_6871_9117# 0.311f
C806 counter\[8\] net6 0.889f
C807 a_4885_7125# _006_ 0.188f
C808 net9 _026_ 0.489f
C809 VPWR a_1547_10004# 0.284f
C810 net9 clknet_1_0__leaf_clk 0.147f
C811 net14 a_4351_2773# 0.439f
C812 _068_ counter\[4\] 1.2f
C813 _056_ clknet_1_1__leaf_clk 0.157f
C814 VPWR a_7619_8916# 0.2f
C815 VPWR a_7090_4765# 0.254f
C816 a_3061_9411# a_2961_9295# 0.168f
C817 net1 net10 0.153f
C818 net14 ones[9] 0.113f
C819 _053_ _025_ 0.407f
C820 _002_ _004_ 0.401f
C821 _063_ _025_ 0.646f
C822 net4 net5 1.06f
C823 _039_ net3 0.184f
C824 net9 counter\[7\] 0.121f
C825 _086_ counter\[0\] 0.397f
C826 VPWR a_9043_3561# 0.202f
C827 net6 _050_ 0.115f
C828 _058_ net7 0.365f
C829 net9 a_5126_5487# 0.166f
C830 a_1925_2473# _093_ 0.108f
C831 _052_ _022_ 0.219f
C832 ones[7] net4 0.451f
C833 a_5639_3311# a_5805_3311# 0.965f
C834 VPWR a_8355_5175# 0.366f
C835 a_4351_2773# a_4958_2741# 0.136f
C836 _037_ a_2419_4221# 0.111f
C837 _043_ _040_ 0.273f
C838 VPWR a_5805_3311# 0.281f
C839 _068_ _055_ 0.181f
C840 a_3243_11293# _060_ 0.217f
C841 net13 net4 0.444f
C842 net13 _042_ 0.117f
C843 VPWR ready 0.219f
C844 VPWR a_2736_9001# 0.164f
C845 net3 _087_ 0.158f
C846 _086_ _050_ 0.157f
C847 counter\[1\] _057_ 0.185f
C848 VPWR _018_ 0.448f
C849 _092_ counter\[0\] 0.295f
C850 VPWR a_8834_8329# 0.31f
C851 net1 counter\[0\] 0.298f
C852 a_8827_8425# a_8834_8329# 0.97f
C853 _088_ a_5177_2487# 0.219f
C854 a_4227_9513# a_4434_9572# 0.26f
C855 net5 ones[3] 0.102f
C856 _057_ counter\[3\] 0.268f
C857 _001_ _060_ 0.115f
C858 a_6987_5161# a_6994_5065# 0.962f
C859 counter\[9\] _040_ 0.793f
C860 a_4234_9417# _028_ 0.113f
C861 _015_ net3 0.327f
C862 _019_ clknet_1_1__leaf_clk 0.212f
C863 a_2603_4405# _031_ 0.117f
C864 VPWR _027_ 1.27f
C865 net4 _039_ 0.372f
C866 VPWR a_4053_6005# 1.21f
C867 VPWR a_7423_10205# 0.179f
C868 VPWR _041_ 0.811f
C869 _048_ _075_ 0.245f
C870 net9 _058_ 0.114f
C871 _090_ _087_ 0.915f
C872 net6 a_7019_2773# 0.424f
C873 counter\[1\] a_1475_5461# 0.128f
C874 _032_ _078_ 2.17f
C875 VPWR a_7527_4087# 0.191f
C876 _072_ counter\[2\] 0.126f
C877 clk VPWR 0.989f
C878 counter\[1\] net13 0.594f
C879 _058_ _054_ 0.368f
C880 clk _070_ 0.187f
C881 VPWR _046_ 1.12f
C882 _091_ _086_ 0.454f
C883 net6 a_9655_9813# 0.248f
C884 a_1761_2767# _007_ 0.121f
C885 net14 _028_ 0.194f
C886 _014_ _083_ 0.142f
C887 VPWR a_1867_9295# 0.27f
C888 _086_ _068_ 0.382f
C889 _073_ net9 0.137f
C890 a_8447_8439# counter\[5\] 0.105f
C891 _041_ net10 0.988f
C892 net3 a_2051_3855# 0.114f
C893 a_1547_10004# _082_ 0.193f
C894 _012_ clk 0.737f
C895 VPWR a_2419_4221# 0.396f
C896 VPWR a_8079_9527# 0.213f
C897 a_7619_8916# _089_ 0.185f
C898 a_8143_6005# counter\[2\] 0.109f
C899 _069_ _007_ 2.05f
C900 a_8022_7119# _037_ 0.13f
C901 _073_ _056_ 0.89f
C902 net6 ones[2] 0.11f
C903 VPWR a_4455_7663# 0.181f
C904 _025_ counter\[6\] 0.248f
C905 _083_ net6 0.106f
C906 _062_ _041_ 0.145f
C907 net10 a_2419_4221# 0.165f
C908 ones[10] _020_ 0.447f
C909 _016_ net14 0.246f
C910 a_8951_10927# a_9390_11293# 0.26f
C911 _090_ _038_ 0.466f
C912 _091_ _092_ 0.134f
C913 _046_ _059_ 0.116f
C914 net7 net11 0.752f
C915 VPWR net12 1.58f
C916 a_6651_4399# _002_ 0.382f
C917 counter\[1\] a_2472_10901# 0.111f
C918 VPWR a_7194_5220# 0.249f
C919 _091_ net1 0.286f
C920 _068_ _092_ 0.981f
C921 _025_ clknet_1_1__leaf_clk 0.115f
C922 _065_ a_4053_6005# 0.137f
C923 VPWR a_3943_9527# 0.168f
C924 a_4338_8751# counter\[4\] 0.102f
C925 _093_ _028_ 0.128f
C926 a_2472_10901# counter\[3\] 0.131f
C927 _060_ clknet_1_1__leaf_clk 0.639f
C928 a_3932_2883# _023_ 0.105f
C929 clknet_1_0__leaf_clk _023_ 0.537f
C930 _092_ _044_ 0.942f
C931 _005_ _060_ 0.161f
C932 _090_ _013_ 0.204f
C933 ones[9] net3 0.225f
C934 counter\[10\] _076_ 0.591f
C935 VPWR _075_ 0.266f
C936 net12 _036_ 0.633f
C937 counter\[1\] _087_ 1.08f
C938 VPWR a_4885_7125# 0.303f
C939 _026_ _025_ 0.378f
C940 _083_ _086_ 0.754f
C941 _014_ a_6361_8751# 0.115f
C942 _039_ net2 0.173f
C943 _090_ _084_ 0.117f
C944 net4 a_8307_10383# 0.189f
C945 counter\[7\] _023_ 0.156f
C946 a_1407_2773# a_2014_2741# 0.141f
C947 _086_ _043_ 0.158f
C948 VPWR _007_ 0.84f
C949 net1 a_9655_9813# 0.178f
C950 _026_ _060_ 0.437f
C951 ones[5] ones[4] 0.112f
C952 VPWR a_9919_8903# 0.219f
C953 _053_ _055_ 0.275f
C954 net13 _052_ 0.217f
C955 clknet_1_0__leaf_clk _060_ 0.215f
C956 a_8355_5175# a_8451_5175# 0.311f
C957 VPWR a_3943_5175# 0.195f
C958 _000_ _085_ 0.102f
C959 net12 _059_ 0.811f
C960 counter\[8\] a_7527_4087# 0.175f
C961 _002_ counter\[5\] 0.596f
C962 VPWR a_7111_10383# 0.303f
C963 VPWR _022_ 1.49f
C964 VPWR a_8022_7119# 1.28f
C965 counter\[10\] _031_ 0.133f
C966 _046_ _033_ 0.162f
C967 _002_ clknet_1_1__leaf_clk 0.435f
C968 _031_ _023_ 0.197f
C969 _009_ net7 0.359f
C970 a_8583_6397# counter\[5\] 0.217f
C971 a_4885_7125# a_4719_7125# 0.966f
C972 _086_ counter\[9\] 0.351f
C973 net1 ones[2] 0.132f
C974 net12 _080_ 0.669f
C975 a_8583_6397# counter\[6\] 0.109f
C976 _025_ counter\[2\] 0.192f
C977 _036_ _022_ 0.105f
C978 _071_ _042_ 1.19f
C979 _056_ a_1665_10383# 0.152f
C980 _067_ _038_ 0.162f
C981 a_6651_4399# a_6817_4399# 0.962f
C982 net14 a_5383_2741# 0.162f
C983 _046_ _050_ 0.288f
C984 a_6803_9513# clknet_1_1__leaf_clk 0.283f
C985 a_7975_6031# a_7277_6037# 0.192f
C986 a_8742_5065# VPWR 0.278f
C987 _001_ _055_ 0.382f
C988 _004_ a_6987_5161# 0.161f
C989 VPWR a_8963_8585# 0.188f
C990 a_7363_5461# VPWR 0.45f
C991 VPWR _000_ 0.515f
C992 VPWR a_4434_6549# 0.242f
C993 _070_ _000_ 0.522f
C994 a_8951_10927# net14 0.401f
C995 a_8827_8425# a_8963_8585# 0.141f
C996 a_4234_9417# a_4363_9673# 0.114f
C997 a_4873_7663# _004_ 0.115f
C998 a_2063_5487# VPWR 0.216f
C999 a_2736_9001# _044_ 0.106f
C1000 _008_ a_7895_8916# 0.109f
C1001 VPWR a_6423_9527# 0.384f
C1002 VPWR a_8815_9527# 0.204f
C1003 net9 net7 0.168f
C1004 _091_ _027_ 1.43f
C1005 counter\[1\] a_4043_10901# 0.202f
C1006 VPWR a_7185_2773# 0.308f
C1007 net11 _029_ 0.221f
C1008 net4 _030_ 0.151f
C1009 _066_ _026_ 0.466f
C1010 _091_ _041_ 0.154f
C1011 a_9919_8439# _063_ 0.204f
C1012 a_4517_2773# a_5215_2767# 0.192f
C1013 VPWR a_7111_6037# 0.452f
C1014 a_4434_5220# VPWR 0.247f
C1015 _041_ _068_ 0.297f
C1016 _061_ net3 1.66f
C1017 a_3775_9527# a_3943_9527# 0.311f
C1018 VPWR a_9209_10389# 0.278f
C1019 net12 _082_ 0.151f
C1020 counter\[5\] counter\[4\] 1.44f
C1021 a_7847_10383# _051_ 0.186f
C1022 _080_ _022_ 0.373f
C1023 _078_ _028_ 0.288f
C1024 net12 _050_ 0.2f
C1025 _084_ counter\[3\] 0.1f
C1026 a_1407_8213# a_2014_8181# 0.141f
C1027 _019_ clknet_0_clk 0.16f
C1028 VPWR a_3847_6727# 0.393f
C1029 a_7822_5761# a_7815_5461# 0.965f
C1030 a_5411_7815# _075_ 0.22f
C1031 _068_ a_7527_4087# 0.196f
C1032 clk _068_ 0.209f
C1033 counter\[4\] clknet_1_1__leaf_clk 0.11f
C1034 net13 a_8583_10927# 0.186f
C1035 _071_ counter\[3\] 0.595f
C1036 clknet_1_1__leaf_clk a_6817_4399# 0.332f
C1037 VPWR a_2736_5059# 0.172f
C1038 a_4319_7637# counter\[4\] 0.309f
C1039 a_4627_8320# _028_ 0.213f
C1040 VPWR a_10239_7663# 0.287f
C1041 a_1925_2473# net2 0.191f
C1042 _073_ _060_ 0.115f
C1043 _066_ counter\[2\] 0.132f
C1044 VPWR a_2439_2741# 0.432f
C1045 _077_ _078_ 0.178f
C1046 _026_ counter\[4\] 1.56f
C1047 clknet_1_0__leaf_clk counter\[4\] 0.2f
C1048 _014_ counter\[5\] 0.244f
C1049 VPWR _057_ 0.742f
C1050 a_8079_9527# a_8352_9527# 0.168f
C1051 VPWR a_6009_10089# 0.227f
C1052 counter\[6\] _055_ 0.422f
C1053 a_6173_8751# _042_ 0.182f
C1054 net10 a_10239_7663# 0.226f
C1055 a_7363_5461# counter\[0\] 0.126f
C1056 VPWR net5 2.61f
C1057 a_3847_5175# a_3943_5175# 0.311f
C1058 _070_ net5 0.343f
C1059 counter\[7\] counter\[4\] 0.217f
C1060 _041_ _083_ 0.144f
C1061 clknet_1_0__leaf_clk _049_ 0.117f
C1062 VPWR a_9135_5737# 0.205f
C1063 net9 _054_ 0.127f
C1064 _014_ clknet_1_1__leaf_clk 0.183f
C1065 _055_ clknet_1_1__leaf_clk 0.157f
C1066 a_5077_2269# a_5177_2487# 0.168f
C1067 _061_ _042_ 0.289f
C1068 _018_ _074_ 0.157f
C1069 _012_ net5 0.241f
C1070 _057_ _036_ 0.38f
C1071 VPWR ones[7] 0.416f
C1072 net4 _028_ 0.189f
C1073 counter\[8\] a_6423_9527# 0.13f
C1074 _057_ net10 0.236f
C1075 a_4326_7937# VPWR 0.282f
C1076 _067_ net8 0.172f
C1077 net9 _029_ 0.117f
C1078 VPWR a_5158_7119# 0.247f
C1079 VPWR a_1475_5461# 0.471f
C1080 clk _043_ 0.101f
C1081 _091_ _007_ 0.225f
C1082 a_8307_10927# ready 0.111f
C1083 a_5779_5175# _037_ 0.222f
C1084 _093_ net3 0.174f
C1085 clknet_1_1__leaf_clk _017_ 0.185f
C1086 net13 VPWR 2.82f
C1087 a_2603_9839# net3 0.146f
C1088 _068_ _007_ 0.207f
C1089 a_7111_6037# _033_ 0.43f
C1090 VPWR a_4234_5065# 0.295f
C1091 _079_ _075_ 0.14f
C1092 VPWR a_10075_10357# 0.392f
C1093 _012_ net13 0.16f
C1094 _062_ _057_ 0.452f
C1095 counter\[7\] _055_ 0.152f
C1096 net14 net4 0.126f
C1097 a_1407_8213# clknet_1_0__leaf_clk 0.277f
C1098 counter\[10\] net11 0.25f
C1099 counter\[1\] _061_ 0.192f
C1100 _026_ net6 0.268f
C1101 net13 _036_ 1.25f
C1102 _057_ _080_ 0.748f
C1103 a_8742_5065# a_8451_5175# 0.189f
C1104 net11 _023_ 0.522f
C1105 clknet_1_0__leaf_clk net6 0.48f
C1106 _081_ _037_ 0.105f
C1107 net13 net10 0.251f
C1108 net8 net2 0.123f
C1109 VPWR _039_ 1.78f
C1110 a_5158_7119# a_4719_7125# 0.273f
C1111 _061_ counter\[3\] 0.13f
C1112 _025_ net11 0.564f
C1113 _056_ _072_ 0.409f
C1114 net12 _043_ 0.361f
C1115 a_6651_4399# a_7090_4765# 0.26f
C1116 a_10100_7351# a_9827_7351# 0.168f
C1117 net13 _059_ 0.143f
C1118 _038_ _037_ 0.272f
C1119 a_8735_5161# a_8742_5065# 0.966f
C1120 a_2839_7351# VPWR 0.211f
C1121 a_8871_5321# VPWR 0.175f
C1122 net2 a_7431_3285# 0.201f
C1123 _057_ counter\[8\] 0.243f
C1124 VPWR a_2472_10901# 0.155f
C1125 VPWR a_6377_5737# 0.195f
C1126 _002_ a_6099_4399# 0.108f
C1127 VPWR a_9117_10927# 0.292f
C1128 _036_ _039_ 0.36f
C1129 a_7822_5761# VPWR 0.298f
C1130 VPWR _003_ 0.351f
C1131 counter\[8\] net5 0.375f
C1132 _008_ a_6803_9513# 0.137f
C1133 a_6939_9673# a_6810_9417# 0.119f
C1134 a_9034_8484# a_8963_8585# 0.24f
C1135 clknet_1_0__leaf_clk _086_ 0.376f
C1136 a_10239_9295# ones[7] 0.11f
C1137 _039_ net10 0.834f
C1138 _077_ _067_ 0.534f
C1139 VPWR a_7458_2767# 0.242f
C1140 _093_ _042_ 0.122f
C1141 a_1407_7119# net2 0.206f
C1142 VPWR _087_ 1.56f
C1143 net13 _080_ 0.617f
C1144 ones[1] a_10239_2223# 0.119f
C1145 _004_ _075_ 0.118f
C1146 clknet_0_clk _066_ 0.138f
C1147 _022_ _045_ 0.171f
C1148 a_2134_5461# a_2063_5487# 0.24f
C1149 net12 counter\[9\] 0.173f
C1150 _028_ net2 0.667f
C1151 _086_ counter\[7\] 0.434f
C1152 clknet_1_1__leaf_clk a_6987_5161# 0.604f
C1153 a_8742_5065# _021_ 0.236f
C1154 a_5779_5175# VPWR 0.201f
C1155 net7 _060_ 0.331f
C1156 VPWR a_1846_8207# 0.287f
C1157 a_8815_9527# _044_ 0.201f
C1158 a_6007_8751# a_6173_8751# 0.959f
C1159 _088_ _017_ 0.392f
C1160 net13 counter\[0\] 0.285f
C1161 a_7019_2773# a_7185_2773# 0.968f
C1162 net5 _050_ 0.917f
C1163 _058_ _055_ 1.16f
C1164 _027_ _047_ 0.38f
C1165 _062_ _039_ 0.123f
C1166 a_7111_10383# _043_ 0.103f
C1167 VPWR _015_ 0.506f
C1168 _036_ _087_ 0.119f
C1169 VPWR a_4234_6849# 0.268f
C1170 a_7822_5761# a_7951_5487# 0.111f
C1171 net13 counter\[8\] 0.227f
C1172 a_6375_7119# _048_ 0.203f
C1173 net8 _034_ 0.263f
C1174 ones[7] _082_ 0.391f
C1175 _042_ a_9279_8725# 0.114f
C1176 _086_ counter\[2\] 0.168f
C1177 net5 _024_ 0.367f
C1178 net1 a_3932_2883# 0.138f
C1179 net1 clknet_1_0__leaf_clk 0.398f
C1180 VPWR _081_ 0.428f
C1181 ones[4] a_10239_5487# 0.11f
C1182 _073_ _055_ 1.47f
C1183 a_4885_7125# a_5326_7093# 0.111f
C1184 net14 net2 0.355f
C1185 _081_ a_6559_9839# 0.113f
C1186 net8 a_7815_5461# 0.101f
C1187 _001_ clk 1.43f
C1188 _077_ net2 0.424f
C1189 a_8583_10927# ones[9] 0.118f
C1190 _058_ _017_ 0.394f
C1191 VPWR _032_ 1.69f
C1192 _032_ _070_ 0.116f
C1193 net13 _082_ 0.182f
C1194 VPWR a_2957_2999# 0.16f
C1195 _086_ _088_ 0.124f
C1196 net9 counter\[10\] 0.438f
C1197 net13 _050_ 0.664f
C1198 net1 counter\[7\] 0.529f
C1199 VPWR _038_ 1.14f
C1200 _032_ a_1499_6031# 0.181f
C1201 VPWR a_2051_3855# 0.179f
C1202 VPWR a_8307_10383# 0.2f
C1203 a_2472_10901# counter\[0\] 0.125f
C1204 _015_ _059_ 0.17f
C1205 _091_ net5 0.655f
C1206 _068_ net5 0.254f
C1207 a_3677_7497# _013_ 0.115f
C1208 net14 _006_ 0.335f
C1209 _035_ _034_ 0.592f
C1210 net9 _060_ 0.53f
C1211 VPWR _013_ 0.864f
C1212 VPWR a_4043_10901# 0.477f
C1213 a_6546_5487# net8 0.23f
C1214 net1 counter\[2\] 1.01f
C1215 _075_ a_4338_8751# 0.113f
C1216 _058_ _086_ 0.129f
C1217 VPWR a_7277_6037# 0.303f
C1218 a_1925_2473# VPWR 0.204f
C1219 _009_ a_4781_5321# 0.118f
C1220 VPWR _084_ 1.46f
C1221 _018_ clknet_1_1__leaf_clk 0.118f
C1222 net12 _047_ 0.12f
C1223 _093_ net2 1.31f
C1224 net7 _040_ 0.268f
C1225 a_4526_7637# VPWR 0.245f
C1226 net1 _088_ 0.2f
C1227 _005_ a_8834_8329# 0.265f
C1228 ones[6] net4 0.193f
C1229 net11 counter\[4\] 0.176f
C1230 VPWR a_1934_5761# 0.352f
C1231 net5 a_9655_9813# 0.156f
C1232 VPWR a_6939_9673# 0.206f
C1233 VPWR _071_ 1.26f
C1234 _056_ _060_ 0.114f
C1235 net14 _034_ 0.171f
C1236 a_2695_6144# _060_ 0.249f
C1237 a_2473_6549# _049_ 0.154f
C1238 _084_ _036_ 1.28f
C1239 a_6519_9527# a_6810_9417# 0.193f
C1240 VPWR a_6375_7119# 0.274f
C1241 VPWR a_4351_2773# 0.399f
C1242 _084_ net10 1.58f
C1243 a_3179_6031# _084_ 0.104f
C1244 VPWR ones[9] 0.344f
C1245 ones[8] net11 0.144f
C1246 _050_ _087_ 0.846f
C1247 a_6546_5487# _035_ 0.147f
C1248 net8 _085_ 0.165f
C1249 VPWR _030_ 1.89f
C1250 a_5607_11079# _086_ 0.181f
C1251 clknet_1_0__leaf_clk _027_ 0.613f
C1252 _070_ _030_ 2.49f
C1253 net7 a_6817_4399# 0.155f
C1254 _084_ a_6835_3968# 0.232f
C1255 _091_ _039_ 0.215f
C1256 _057_ _043_ 0.148f
C1257 a_4053_6005# clknet_1_0__leaf_clk 1.64f
C1258 _028_ _037_ 0.644f
C1259 net11 _055_ 0.27f
C1260 a_4434_5220# a_4227_5161# 0.26f
C1261 VPWR a_1669_6727# 0.184f
C1262 a_3130_7241# VPWR 0.328f
C1263 a_8735_5161# a_8871_5321# 0.136f
C1264 _082_ _081_ 0.172f
C1265 _093_ _034_ 0.662f
C1266 _084_ _080_ 0.135f
C1267 a_9397_10383# _020_ 0.114f
C1268 VPWR a_9390_11293# 0.235f
C1269 _046_ _026_ 0.537f
C1270 _038_ _033_ 0.109f
C1271 counter\[1\] net3 0.199f
C1272 a_4043_10901# counter\[0\] 0.233f
C1273 _009_ counter\[4\] 1.06f
C1274 _046_ clknet_1_0__leaf_clk 0.321f
C1275 _081_ a_6178_9839# 0.114f
C1276 clk _076_ 0.479f
C1277 _048_ net14 0.112f
C1278 a_7363_5461# a_7531_5461# 0.311f
C1279 _013_ counter\[8\] 0.13f
C1280 counter\[3\] net3 0.112f
C1281 a_2695_6144# _066_ 0.202f
C1282 a_4434_6549# a_4363_6575# 0.24f
C1283 net7 a_10239_4399# 0.195f
C1284 net14 _037_ 0.162f
C1285 _014_ net7 0.104f
C1286 VPWR net8 1.54f
C1287 a_4319_7637# a_4455_7663# 0.136f
C1288 a_4326_7937# _004_ 0.281f
C1289 counter\[9\] net5 0.205f
C1290 _084_ counter\[8\] 0.14f
C1291 net12 clknet_1_1__leaf_clk 0.105f
C1292 net13 _043_ 0.145f
C1293 VPWR a_2271_8207# 0.194f
C1294 VPWR a_7431_3285# 0.204f
C1295 a_7019_2773# a_7458_2767# 0.26f
C1296 a_7185_2773# a_7626_2741# 0.127f
C1297 VPWR a_6173_8751# 0.309f
C1298 net2 net3 0.522f
C1299 net12 _026_ 0.225f
C1300 a_9728_6147# _025_ 0.123f
C1301 VPWR a_1407_10927# 0.365f
C1302 net6 net7 0.149f
C1303 clknet_1_0__leaf_clk net12 0.805f
C1304 _009_ _014_ 0.482f
C1305 VPWR _061_ 0.746f
C1306 a_4035_7637# a_4326_7937# 0.192f
C1307 VPWR a_1407_7119# 0.391f
C1308 a_1669_6727# _080_ 0.107f
C1309 net12 _076_ 0.29f
C1310 a_5326_7093# a_5158_7119# 0.24f
C1311 a_4434_5220# a_4363_5321# 0.24f
C1312 VPWR a_4234_9417# 0.274f
C1313 _015_ a_7019_2773# 0.138f
C1314 a_9427_9295# _028_ 0.214f
C1315 _071_ _082_ 0.129f
C1316 VPWR _028_ 3.22f
C1317 VPWR a_6519_9527# 0.176f
C1318 a_9209_10389# a_9650_10357# 0.127f
C1319 _008_ a_7619_8916# 0.123f
C1320 VPWR _035_ 1.67f
C1321 counter\[1\] net4 0.225f
C1322 VPWR a_9137_7913# 0.243f
C1323 a_5583_7119# a_4885_7125# 0.195f
C1324 a_1407_8213# a_1573_8213# 0.969f
C1325 _091_ a_2051_3855# 0.128f
C1326 a_2743_7351# net6 0.107f
C1327 _075_ _076_ 0.105f
C1328 a_1669_6727# counter\[8\] 0.207f
C1329 VPWR a_9043_10389# 0.395f
C1330 a_8022_7119# clknet_1_1__leaf_clk 1.67f
C1331 _003_ _043_ 0.203f
C1332 _042_ counter\[3\] 0.235f
C1333 a_7039_9019# net7 0.15f
C1334 counter\[10\] _060_ 0.313f
C1335 clknet_1_0__leaf_clk _007_ 0.119f
C1336 net9 _055_ 0.148f
C1337 a_3847_6727# a_3943_6549# 0.311f
C1338 _001_ a_2481_5487# 0.119f
C1339 _016_ a_5639_3311# 0.131f
C1340 a_3130_7241# counter\[8\] 0.245f
C1341 net11 a_7591_10107# 0.142f
C1342 _035_ _036_ 0.116f
C1343 _049_ _029_ 0.485f
C1344 a_4227_5161# a_4234_5065# 0.963f
C1345 a_6078_3677# a_5639_3311# 0.26f
C1346 a_6246_3423# a_5805_3311# 0.111f
C1347 _053_ net13 0.28f
C1348 net14 a_9427_9295# 0.103f
C1349 net12 _031_ 0.145f
C1350 a_6377_5737# _074_ 0.128f
C1351 VPWR net14 4.7f
C1352 net1 net11 0.129f
C1353 _035_ net10 0.192f
C1354 _089_ _030_ 0.113f
C1355 _000_ counter\[5\] 1.04f
C1356 a_4043_10901# _068_ 0.114f
C1357 _025_ _060_ 0.263f
C1358 _077_ VPWR 1.29f
C1359 _016_ VPWR 0.43f
C1360 a_6871_9117# a_6173_8751# 0.192f
C1361 clknet_1_0__leaf_clk _022_ 0.224f
C1362 VPWR a_6078_3677# 0.249f
C1363 _003_ _074_ 0.878f
C1364 a_4903_4399# _078_ 0.203f
C1365 a_8742_5065# clknet_1_1__leaf_clk 0.29f
C1366 ones[10] ready 0.166f
C1367 _012_ net14 0.133f
C1368 _084_ _068_ 0.957f
C1369 _034_ net3 0.487f
C1370 _056_ _055_ 0.388f
C1371 net4 net2 0.418f
C1372 net9 a_5316_5487# 0.117f
C1373 _022_ counter\[7\] 0.344f
C1374 VPWR a_1573_2773# 0.35f
C1375 a_4234_6849# _043_ 0.349f
C1376 _062_ _028_ 0.201f
C1377 _068_ _071_ 0.102f
C1378 net14 net10 0.127f
C1379 net8 _033_ 0.13f
C1380 VPWR a_6375_4399# 0.198f
C1381 _054_ _017_ 0.147f
C1382 _010_ _032_ 1.3f
C1383 a_4781_9673# _011_ 0.119f
C1384 VPWR a_4958_2741# 0.184f
C1385 _032_ _083_ 0.394f
C1386 _080_ _028_ 1.18f
C1387 VPWR a_9827_7351# 0.213f
C1388 counter\[1\] counter\[3\] 1.15f
C1389 a_7111_6037# clknet_1_1__leaf_clk 0.25f
C1390 net14 _059_ 0.355f
C1391 _004_ _081_ 0.235f
C1392 a_2439_2741# a_2271_2767# 0.311f
C1393 a_9209_10389# clknet_1_1__leaf_clk 0.181f
C1394 _016_ _059_ 0.732f
C1395 net8 _050_ 0.184f
C1396 _014_ _072_ 0.83f
C1397 a_8735_5161# _030_ 0.437f
C1398 VPWR _093_ 1.7f
C1399 VPWR a_2603_9839# 0.404f
C1400 VPWR a_2375_10615# 0.207f
C1401 _062_ net14 0.12f
C1402 net4 _052_ 0.369f
C1403 counter\[8\] _028_ 0.12f
C1404 a_4053_6005# clknet_0_clk 0.343f
C1405 _012_ _093_ 0.64f
C1406 a_5805_3311# net11 0.104f
C1407 _035_ counter\[8\] 0.441f
C1408 VPWR a_3247_6575# 0.24f
C1409 a_4363_5321# a_4234_5065# 0.119f
C1410 net14 _080_ 1.03f
C1411 counter\[10\] _040_ 0.516f
C1412 a_2736_9001# net11 0.174f
C1413 _010_ _084_ 0.241f
C1414 VPWR a_1499_10383# 0.23f
C1415 _061_ _082_ 1.86f
C1416 a_8942_5220# a_8871_5321# 0.24f
C1417 a_9209_10389# a_9907_10383# 0.194f
C1418 _040_ _023_ 0.106f
C1419 _061_ _089_ 0.129f
C1420 VPWR a_7550_6031# 0.255f
C1421 counter\[9\] a_2957_2999# 0.184f
C1422 _066_ _060_ 0.416f
C1423 clk clknet_0_clk 0.231f
C1424 _037_ net3 0.531f
C1425 VPWR a_5383_2741# 0.434f
C1426 VPWR a_9279_8725# 0.417f
C1427 net14 counter\[0\] 0.178f
C1428 _082_ _028_ 0.282f
C1429 _000_ counter\[2\] 0.166f
C1430 counter\[9\] _038_ 0.159f
C1431 _009_ a_7619_8916# 0.111f
C1432 _050_ _028_ 0.412f
C1433 net5 counter\[6\] 0.355f
C1434 _026_ a_2736_5059# 0.166f
C1435 a_7531_5461# a_7822_5761# 0.195f
C1436 _035_ _089_ 0.489f
C1437 _027_ net11 0.205f
C1438 _040_ _060_ 0.109f
C1439 a_8951_10927# VPWR 0.457f
C1440 counter\[1\] _006_ 0.372f
C1441 _084_ _074_ 0.184f
C1442 VPWR a_10239_3311# 0.281f
C1443 a_7626_2741# a_7458_2767# 0.24f
C1444 _057_ clknet_1_0__leaf_clk 0.109f
C1445 VPWR a_10239_6575# 0.275f
C1446 _026_ net5 0.304f
C1447 clknet_1_0__leaf_clk net5 0.962f
C1448 net7 _027_ 0.312f
C1449 VPWR a_3970_9839# 0.206f
C1450 a_4434_6549# a_4227_6549# 0.26f
C1451 a_4363_6575# a_4234_6849# 0.119f
C1452 a_1669_6727# _083_ 0.138f
C1453 a_4326_7937# a_4319_7637# 0.967f
C1454 _061_ _068_ 0.203f
C1455 counter\[9\] _071_ 0.578f
C1456 a_3061_9411# _029_ 0.114f
C1457 _093_ counter\[0\] 0.108f
C1458 VPWR a_4363_9673# 0.174f
C1459 _092_ _011_ 0.216f
C1460 _091_ _028_ 0.699f
C1461 net13 clknet_1_1__leaf_clk 0.295f
C1462 a_2014_8181# a_1846_8207# 0.24f
C1463 a_1475_5461# a_1643_5461# 0.311f
C1464 VPWR a_4993_3855# 0.19f
C1465 VPWR a_9983_11195# 0.454f
C1466 a_4326_7937# _026_ 0.212f
C1467 _061_ _044_ 0.512f
C1468 _042_ _037_ 0.209f
C1469 VPWR ones[6] 0.293f
C1470 _052_ net2 0.101f
C1471 a_9827_7351# _082_ 0.126f
C1472 a_1499_10383# counter\[0\] 0.288f
C1473 _028_ _044_ 0.506f
C1474 net13 _026_ 0.207f
C1475 VPWR _078_ 0.64f
C1476 VPWR a_2691_6825# 0.265f
C1477 VPWR net3 4.51f
C1478 _079_ _028_ 0.328f
C1479 net13 clknet_1_0__leaf_clk 0.265f
C1480 _010_ net8 0.499f
C1481 _070_ net3 0.344f
C1482 _035_ _044_ 0.143f
C1483 a_2971_3311# _015_ 0.109f
C1484 a_3943_6549# a_4234_6849# 0.192f
C1485 VPWR a_5915_5487# 0.189f
C1486 _025_ _055_ 0.153f
C1487 net7 a_2419_4221# 0.138f
C1488 _012_ _078_ 0.273f
C1489 net12 net11 0.361f
C1490 _091_ net14 0.101f
C1491 _012_ net3 0.412f
C1492 net14 _068_ 0.131f
C1493 _014_ _060_ 0.527f
C1494 a_4517_2773# _022_ 0.178f
C1495 a_10075_10357# a_9907_10383# 0.311f
C1496 _002_ counter\[4\] 0.219f
C1497 VPWR a_9963_2223# 0.27f
C1498 VPWR a_6503_3677# 0.197f
C1499 VPWR a_4627_8320# 0.258f
C1500 _036_ net3 0.219f
C1501 a_8022_7119# clknet_0_clk 0.314f
C1502 VPWR a_3063_11293# 0.203f
C1503 net6 _023_ 0.127f
C1504 a_9117_10927# clknet_1_1__leaf_clk 0.203f
C1505 _026_ _039_ 0.177f
C1506 net8 _074_ 0.179f
C1507 _077_ _079_ 0.134f
C1508 _025_ net6 0.402f
C1509 _001_ _084_ 0.238f
C1510 a_2439_8181# net5 0.127f
C1511 a_8583_6397# counter\[4\] 0.143f
C1512 net12 net7 0.117f
C1513 _090_ VPWR 0.507f
C1514 _059_ net3 0.285f
C1515 _060_ _017_ 0.914f
C1516 _058_ _057_ 0.161f
C1517 net8 counter\[9\] 0.248f
C1518 net6 _060_ 0.203f
C1519 a_2795_4649# VPWR 0.126f
C1520 a_7718_6005# a_7111_6037# 0.136f
C1521 _001_ a_1934_5761# 0.244f
C1522 a_4864_3829# _023_ 0.152f
C1523 a_2063_5487# a_1927_5461# 0.141f
C1524 _043_ _028_ 0.435f
C1525 _003_ clknet_1_0__leaf_clk 0.114f
C1526 net4 a_5639_3311# 0.45f
C1527 VPWR a_10100_7351# 0.184f
C1528 clk net9 0.11f
C1529 counter\[1\] _069_ 0.189f
C1530 _091_ _093_ 0.123f
C1531 _027_ _029_ 1.28f
C1532 _015_ clknet_1_1__leaf_clk 0.148f
C1533 VPWR net4 6f
C1534 VPWR _042_ 2.74f
C1535 _090_ a_3179_6031# 0.147f
C1536 clknet_1_0__leaf_clk _087_ 0.391f
C1537 _080_ net3 0.109f
C1538 a_6446_9117# a_6007_8751# 0.26f
C1539 _049_ _040_ 0.197f
C1540 _009_ net12 0.119f
C1541 clk _054_ 0.114f
C1542 _074_ _028_ 0.18f
C1543 _053_ net8 0.263f
C1544 _081_ clknet_1_1__leaf_clk 0.324f
C1545 a_1867_9295# _054_ 0.191f
C1546 a_9919_8439# _060_ 0.188f
C1547 counter\[0\] net3 0.111f
C1548 _013_ a_4767_5652# 0.107f
C1549 net4 _036_ 0.25f
C1550 net7 _022_ 1.19f
C1551 a_2472_10901# counter\[2\] 0.141f
C1552 counter\[8\] net3 0.106f
C1553 VPWR a_7975_6031# 0.174f
C1554 _009_ _075_ 0.277f
C1555 a_9117_10927# a_9558_11039# 0.125f
C1556 VPWR a_6375_2775# 0.292f
C1557 _004_ net14 0.194f
C1558 _003_ counter\[2\] 0.293f
C1559 _000_ a_8215_8751# 0.109f
C1560 a_3775_9527# net3 0.154f
C1561 ones[6] _082_ 0.122f
C1562 counter\[0\] a_3063_11293# 0.245f
C1563 _065_ _090_ 0.178f
C1564 counter\[2\] _087_ 0.156f
C1565 _048_ _006_ 0.479f
C1566 VPWR a_6725_9839# 0.292f
C1567 _082_ net3 0.429f
C1568 VPWR _067_ 1.45f
C1569 counter\[1\] VPWR 2.43f
C1570 a_6725_9839# a_6559_9839# 0.966f
C1571 VPWR ones[3] 0.308f
C1572 VPWR a_8051_2741# 0.409f
C1573 clknet_1_0__leaf_clk _038_ 0.616f
C1574 _063_ _028_ 0.201f
C1575 _001_ net8 1.7f
C1576 _000_ net7 0.256f
C1577 a_10100_7351# _080_ 0.124f
C1578 VPWR counter\[3\] 0.904f
C1579 _071_ counter\[6\] 0.142f
C1580 _005_ _084_ 0.314f
C1581 a_9043_10389# a_9482_10383# 0.26f
C1582 _059_ a_6375_2775# 0.175f
C1583 _067_ _036_ 0.271f
C1584 net3 _024_ 0.181f
C1585 net12 _029_ 0.254f
C1586 a_8307_10927# net14 0.223f
C1587 _003_ a_4227_6549# 0.1f
C1588 _013_ clknet_1_0__leaf_clk 0.659f
C1589 _055_ _051_ 0.107f
C1590 a_4319_7637# a_4526_7637# 0.26f
C1591 _034_ _037_ 0.17f
C1592 _067_ a_3179_6031# 0.178f
C1593 counter\[1\] net10 0.273f
C1594 counter\[2\] _081_ 0.423f
C1595 _038_ a_5126_5487# 0.11f
C1596 net4 counter\[0\] 0.131f
C1597 _042_ counter\[0\] 0.134f
C1598 a_6803_9513# a_7010_9572# 0.273f
C1599 _014_ _049_ 1.06f
C1600 _084_ _026_ 0.105f
C1601 _064_ net8 0.159f
C1602 VPWR a_7469_10703# 0.193f
C1603 a_1643_5461# a_1934_5761# 0.197f
C1604 a_9427_9295# net2 0.113f
C1605 counter\[8\] _042_ 0.285f
C1606 VPWR net2 3.01f
C1607 ones[9] clknet_1_1__leaf_clk 0.132f
C1608 _086_ _040_ 0.126f
C1609 VPWR a_8543_8439# 0.21f
C1610 net13 _008_ 0.222f
C1611 _017_ a_6817_4399# 0.174f
C1612 a_5805_3311# _023_ 0.268f
C1613 _091_ net3 1.63f
C1614 _047_ _028_ 0.262f
C1615 _030_ clknet_1_1__leaf_clk 0.346f
C1616 a_1489_4943# VPWR 0.171f
C1617 _062_ counter\[1\] 0.216f
C1618 _088_ a_2957_2999# 0.125f
C1619 a_4234_6849# a_4227_6549# 0.962f
C1620 clknet_1_0__leaf_clk a_4351_2773# 0.334f
C1621 net7 a_2736_5059# 0.18f
C1622 _068_ a_5915_5487# 0.227f
C1623 _073_ _087_ 0.255f
C1624 net5 net11 0.594f
C1625 net6 _049_ 0.481f
C1626 net4 _082_ 0.726f
C1627 a_3130_7241# a_3259_7497# 0.119f
C1628 a_3123_7337# _013_ 0.123f
C1629 _065_ _067_ 0.432f
C1630 a_3247_6575# counter\[9\] 0.234f
C1631 net4 _050_ 0.161f
C1632 VPWR a_7515_4765# 0.187f
C1633 a_4043_10901# counter\[2\] 0.157f
C1634 _065_ counter\[1\] 0.732f
C1635 net4 _089_ 0.556f
C1636 VPWR a_6007_8751# 0.44f
C1637 ones[2] a_10239_3311# 0.11f
C1638 _042_ _089_ 0.297f
C1639 net9 _000_ 0.269f
C1640 _026_ _030_ 0.112f
C1641 VPWR _006_ 0.382f
C1642 _072_ _007_ 2.42f
C1643 _080_ counter\[3\] 0.209f
C1644 VPWR a_5722_6575# 1.23f
C1645 _001_ net14 0.105f
C1646 counter\[1\] counter\[0\] 1.69f
C1647 VPWR _052_ 1.69f
C1648 a_2327_9295# _018_ 0.109f
C1649 net8 counter\[5\] 0.465f
C1650 _032_ _058_ 0.197f
C1651 _019_ net12 0.952f
C1652 a_9043_10389# a_9650_10357# 0.136f
C1653 net13 a_2473_6549# 0.166f
C1654 a_5607_11079# _087_ 0.116f
C1655 _048_ _037_ 0.113f
C1656 net5 net7 0.206f
C1657 _012_ _052_ 1.21f
C1658 _020_ a_9209_10389# 0.18f
C1659 _071_ counter\[2\] 0.176f
C1660 counter\[0\] counter\[3\] 0.758f
C1661 net13 net11 0.153f
C1662 a_10011_5175# _030_ 0.107f
C1663 _010_ a_7541_5321# 0.125f
C1664 net8 clknet_1_1__leaf_clk 0.182f
C1665 _027_ _060_ 0.519f
C1666 a_4903_4399# VPWR 0.247f
C1667 VPWR _034_ 1.52f
C1668 _070_ _034_ 0.108f
C1669 _021_ a_9289_5321# 0.119f
C1670 _003_ clknet_0_clk 0.186f
C1671 VPWR a_9411_2767# 0.259f
C1672 counter\[1\] _082_ 0.114f
C1673 VPWR a_7815_5461# 0.686f
C1674 _083_ net3 0.136f
C1675 _092_ counter\[4\] 1.11f
C1676 _012_ a_9411_2767# 0.112f
C1677 net8 _026_ 0.351f
C1678 a_6173_8751# clknet_1_1__leaf_clk 0.319f
C1679 _031_ _030_ 0.337f
C1680 a_9963_9295# ones[8] 0.114f
C1681 counter\[5\] _028_ 1.38f
C1682 net13 net7 0.128f
C1683 net11 _039_ 0.167f
C1684 counter\[6\] _028_ 0.248f
C1685 a_6446_9117# VPWR 0.258f
C1686 _042_ _044_ 0.111f
C1687 a_3123_7337# a_3130_7241# 0.97f
C1688 VPWR a_6810_9417# 0.296f
C1689 _028_ clknet_1_1__leaf_clk 0.35f
C1690 net6 a_4864_3829# 0.135f
C1691 _005_ _028_ 0.715f
C1692 _078_ _074_ 0.337f
C1693 a_9558_11039# a_9390_11293# 0.24f
C1694 a_6527_6263# _042_ 0.109f
C1695 a_7123_5321# a_6987_5161# 0.141f
C1696 net12 _023_ 0.524f
C1697 a_7815_5461# a_7951_5487# 0.141f
C1698 _086_ net6 0.911f
C1699 a_6546_5487# VPWR 0.203f
C1700 _082_ net2 0.123f
C1701 clknet_0_clk _081_ 0.348f
C1702 _012_ a_1761_8207# 0.116f
C1703 a_2271_2767# a_1573_2773# 0.195f
C1704 net13 _009_ 0.141f
C1705 a_9043_10389# clknet_1_1__leaf_clk 0.308f
C1706 ones[10] a_8307_10383# 0.109f
C1707 counter\[9\] net3 1.56f
C1708 _089_ net2 1.9f
C1709 net14 counter\[6\] 0.894f
C1710 _026_ _028_ 0.566f
C1711 _077_ counter\[6\] 0.102f
C1712 a_4234_5065# _009_ 0.248f
C1713 clknet_1_0__leaf_clk _028_ 0.129f
C1714 VPWR _048_ 0.712f
C1715 net1 _055_ 0.203f
C1716 VPWR a_6998_10205# 0.259f
C1717 _080_ _034_ 0.44f
C1718 a_6998_10205# a_6559_9839# 0.26f
C1719 net12 _060_ 0.144f
C1720 VPWR a_6703_5175# 0.195f
C1721 VPWR _037_ 1.08f
C1722 counter\[1\] _068_ 0.295f
C1723 net14 clknet_1_1__leaf_clk 0.22f
C1724 a_7277_6037# a_7718_6005# 0.111f
C1725 _077_ clknet_1_1__leaf_clk 0.171f
C1726 VPWR a_8583_10927# 0.189f
C1727 net2 _024_ 0.304f
C1728 _039_ a_4719_3311# 0.114f
C1729 _077_ _005_ 0.109f
C1730 _068_ counter\[3\] 0.12f
C1731 _028_ a_10011_5175# 0.17f
C1732 _015_ net11 0.671f
C1733 _035_ counter\[7\] 0.254f
C1734 a_9275_6263# net8 0.223f
C1735 _041_ _040_ 0.196f
C1736 _028_ a_5126_5487# 0.109f
C1737 _069_ VPWR 1.16f
C1738 _075_ _060_ 0.136f
C1739 net4 _043_ 0.397f
C1740 net14 _026_ 0.672f
C1741 _043_ _042_ 1.63f
C1742 _063_ net3 0.116f
C1743 net1 _017_ 0.211f
C1744 net14 a_3932_2883# 0.189f
C1745 net14 clknet_1_0__leaf_clk 0.407f
C1746 a_2839_7351# a_2743_7351# 0.311f
C1747 net11 _081_ 0.298f
C1748 net1 net6 3.71f
C1749 VPWR a_7258_4511# 0.184f
C1750 _052_ _050_ 0.175f
C1751 _022_ _023_ 0.127f
C1752 ones[5] net14 0.126f
C1753 VPWR _085_ 0.764f
C1754 a_2439_8181# a_2271_8207# 0.311f
C1755 _005_ a_6375_4399# 0.109f
C1756 _077_ _076_ 0.1f
C1757 a_1934_5761# a_1927_5461# 0.975f
C1758 clk _040_ 1.06f
C1759 _091_ net2 0.133f
C1760 _046_ _040_ 0.178f
C1761 _047_ a_3970_9839# 0.115f
C1762 net14 counter\[7\] 0.656f
C1763 ones[10] ones[9] 0.222f
C1764 a_7255_3285# a_7431_3285# 0.185f
C1765 _074_ _042_ 0.642f
C1766 clknet_1_0__leaf_clk a_1573_2773# 0.254f
C1767 _022_ _060_ 0.113f
C1768 _058_ a_7431_3285# 0.102f
C1769 a_1489_4943# _068_ 0.163f
C1770 net7 _081_ 0.111f
C1771 a_8815_9527# a_9088_9527# 0.168f
C1772 VPWR a_8079_5162# 0.186f
C1773 a_4351_2773# a_4517_2773# 0.96f
C1774 net10 _085_ 0.418f
C1775 _010_ _067_ 0.601f
C1776 VPWR a_3939_7815# 0.394f
C1777 ones[3] ones[2] 0.112f
C1778 a_6375_4399# _076_ 0.191f
C1779 _066_ net12 0.181f
C1780 _032_ net7 0.584f
C1781 VPWR a_5639_3311# 0.444f
C1782 clk counter\[4\] 0.152f
C1783 a_3243_11293# a_3063_11293# 0.185f
C1784 counter\[1\] _043_ 0.386f
C1785 _046_ counter\[4\] 0.291f
C1786 a_6835_3968# _085_ 0.104f
C1787 VPWR a_9427_9295# 0.349f
C1788 VPWR _070_ 0.844f
C1789 VPWR a_6559_9839# 0.421f
C1790 net12 _040_ 0.625f
C1791 counter\[1\] _004_ 0.101f
C1792 VPWR a_8827_8425# 0.543f
C1793 a_6007_8751# _044_ 0.442f
C1794 _012_ VPWR 2.04f
C1795 _000_ a_8369_5487# 0.137f
C1796 a_4227_9513# a_4234_9417# 0.969f
C1797 VPWR a_1499_6031# 0.233f
C1798 a_4627_8320# _047_ 0.217f
C1799 a_5077_2269# _087_ 0.12f
C1800 a_6703_5175# a_6994_5065# 0.195f
C1801 a_8951_10927# clknet_1_1__leaf_clk 0.305f
C1802 VPWR a_2961_9295# 0.171f
C1803 net1 _092_ 0.119f
C1804 VPWR _036_ 1.49f
C1805 _069_ counter\[0\] 1.77f
C1806 _067_ counter\[9\] 0.209f
C1807 _026_ a_9279_8725# 0.167f
C1808 _068_ _034_ 0.247f
C1809 VPWR net10 2.14f
C1810 counter\[1\] counter\[9\] 0.944f
C1811 _084_ net7 0.307f
C1812 VPWR a_3179_6031# 0.44f
C1813 a_4351_2773# a_4790_2767# 0.26f
C1814 _056_ _087_ 0.587f
C1815 a_1489_4943# a_1589_5059# 0.168f
C1816 VPWR a_7951_5487# 0.184f
C1817 _077_ _058_ 0.182f
C1818 counter\[9\] counter\[3\] 1.55f
C1819 _019_ net13 0.556f
C1820 VPWR _059_ 0.912f
C1821 _016_ a_5993_3311# 0.115f
C1822 _029_ _087_ 1.11f
C1823 VPWR a_4719_7125# 0.693f
C1824 _070_ _059_ 0.205f
C1825 a_8022_7119# _066_ 0.205f
C1826 VPWR a_6835_3968# 0.233f
C1827 a_6871_9117# VPWR 0.215f
C1828 _062_ VPWR 3.28f
C1829 net12 _049_ 0.116f
C1830 _073_ net14 0.124f
C1831 _069_ _082_ 0.254f
C1832 _074_ net2 0.109f
C1833 counter\[1\] _053_ 0.154f
C1834 _075_ counter\[4\] 0.222f
C1835 VPWR a_1632_3971# 0.179f
C1836 net9 _038_ 0.188f
C1837 _078_ counter\[6\] 0.171f
C1838 VPWR _080_ 2.23f
C1839 _065_ VPWR 1.17f
C1840 counter\[5\] a_5915_5487# 0.25f
C1841 ones[5] a_10239_6575# 0.11f
C1842 net7 _030_ 2.04f
C1843 net5 _023_ 1.85f
C1844 _089_ _085_ 1.47f
C1845 a_7123_5321# a_7194_5220# 0.24f
C1846 _066_ _000_ 0.214f
C1847 a_10239_9295# VPWR 0.219f
C1848 _002_ a_7111_6037# 0.117f
C1849 VPWR counter\[0\] 5.73f
C1850 clknet_1_1__leaf_clk net3 0.152f
C1851 _062_ net10 0.208f
C1852 _005_ _078_ 0.918f
C1853 net12 _055_ 0.328f
C1854 VPWR a_9306_7663# 0.221f
C1855 net8 net11 0.191f
C1856 a_8951_10927# a_9558_11039# 0.138f
C1857 _019_ a_9117_10927# 0.18f
C1858 VPWR counter\[8\] 4.75f
C1859 net5 _060_ 0.346f
C1860 VPWR a_6994_5065# 0.317f
C1861 _068_ _037_ 0.667f
C1862 _080_ net10 0.207f
C1863 _038_ _029_ 0.286f
C1864 _053_ a_7469_10703# 0.138f
C1865 net1 ready 0.174f
C1866 net14 ones[10] 0.276f
C1867 _018_ _092_ 0.21f
C1868 a_6246_3423# a_6078_3677# 0.24f
C1869 _052_ _074_ 0.376f
C1870 _043_ _034_ 1.41f
C1871 _012_ counter\[8\] 0.239f
C1872 ones[5] ones[6] 0.112f
C1873 VPWR _033_ 2.49f
C1874 VPWR a_5411_7815# 0.197f
C1875 VPWR a_3775_9527# 0.429f
C1876 _026_ net3 0.212f
C1877 _014_ _075_ 0.162f
C1878 clknet_1_0__leaf_clk net3 0.55f
C1879 _022_ _049_ 0.177f
C1880 _073_ _093_ 0.109f
C1881 counter\[0\] net10 0.398f
C1882 a_7883_2767# a_7185_2773# 0.194f
C1883 VPWR a_4169_9001# 0.268f
C1884 net12 net6 0.48f
C1885 VPWR _082_ 1.66f
C1886 _069_ _068_ 0.193f
C1887 net13 _025_ 0.346f
C1888 net8 net7 0.245f
C1889 VPWR _050_ 1.7f
C1890 a_7423_10205# a_7591_10107# 0.311f
C1891 _055_ a_9919_8903# 0.251f
C1892 VPWR _089_ 0.963f
C1893 _074_ _034_ 1.13f
C1894 _070_ _089_ 0.219f
C1895 _062_ _080_ 0.233f
C1896 _061_ a_8215_8751# 0.188f
C1897 _068_ _085_ 0.307f
C1898 a_1407_2773# a_1573_2773# 0.97f
C1899 net13 _060_ 0.182f
C1900 VPWR a_6178_9839# 0.197f
C1901 net11 _028_ 0.302f
C1902 _041_ net1 0.354f
C1903 VPWR a_3847_5175# 0.418f
C1904 a_9815_11293# a_9117_10927# 0.195f
C1905 VPWR _024_ 0.237f
C1906 _062_ counter\[0\] 1.16f
C1907 _082_ net10 0.126f
C1908 _053_ _052_ 0.115f
C1909 _019_ _081_ 1.1f
C1910 _090_ clknet_1_0__leaf_clk 0.337f
C1911 _050_ net10 1.09f
C1912 _012_ _024_ 0.205f
C1913 _089_ net10 0.341f
C1914 _062_ counter\[8\] 0.646f
C1915 _066_ _057_ 1.73f
C1916 net4 clknet_1_1__leaf_clk 0.135f
C1917 _042_ clknet_1_1__leaf_clk 0.407f
C1918 net8 a_10239_5487# 0.201f
C1919 _080_ counter\[0\] 0.124f
C1920 _065_ counter\[0\] 0.195f
C1921 VPWR a_8451_5175# 0.168f
C1922 a_4517_2773# a_4958_2741# 0.118f
C1923 net7 _028_ 0.701f
C1924 _039_ _060_ 0.169f
C1925 _066_ net5 0.246f
C1926 counter\[8\] _080_ 0.458f
C1927 a_1573_8213# a_2271_8207# 0.195f
C1928 net14 net11 0.36f
C1929 _016_ net11 0.137f
C1930 net6 _022_ 0.128f
C1931 _035_ net7 0.429f
C1932 _043_ _037_ 0.784f
C1933 VPWR _091_ 1.56f
C1934 counter\[10\] _087_ 0.199f
C1935 a_7550_6031# a_7718_6005# 0.24f
C1936 _026_ _042_ 0.195f
C1937 a_9963_9295# net12 0.202f
C1938 a_8735_5161# VPWR 0.394f
C1939 _065_ _033_ 0.184f
C1940 clknet_1_0__leaf_clk net4 0.419f
C1941 VPWR _068_ 3.26f
C1942 net5 _040_ 0.545f
C1943 _070_ _068_ 0.131f
C1944 _064_ net2 1.13f
C1945 ones[5] net4 0.203f
C1946 VPWR a_9034_8484# 0.27f
C1947 _012_ _091_ 0.151f
C1948 net8 net9 0.47f
C1949 a_5779_5175# _023_ 0.205f
C1950 _003_ a_4781_6575# 0.115f
C1951 a_8827_8425# a_9034_8484# 0.273f
C1952 counter\[0\] _033_ 1.11f
C1953 a_4227_9513# a_4363_9673# 0.136f
C1954 a_2134_5461# VPWR 0.272f
C1955 counter\[1\] counter\[6\] 0.332f
C1956 VPWR _044_ 3.25f
C1957 VPWR a_8352_9527# 0.157f
C1958 a_6987_5161# a_7194_5220# 0.26f
C1959 VPWR a_7019_2773# 0.481f
C1960 VPWR _079_ 0.67f
C1961 _077_ net7 1.46f
C1962 _068_ _036_ 0.119f
C1963 _060_ _087_ 0.685f
C1964 a_2795_4649# _031_ 0.132f
C1965 _068_ net10 0.326f
C1966 _077_ a_9544_3561# 0.105f
C1967 counter\[9\] _037_ 0.162f
C1968 a_4958_2741# a_4790_2767# 0.24f
C1969 VPWR a_9655_9813# 0.452f
C1970 VPWR a_6527_6263# 0.204f
C1971 _021_ VPWR 0.174f
C1972 net13 _040_ 0.236f
C1973 counter\[8\] _050_ 0.104f
C1974 _036_ _044_ 0.122f
C1975 a_1665_10383# a_1499_10383# 0.125f
C1976 _068_ _059_ 0.303f
C1977 _019_ a_6375_7119# 0.108f
C1978 _073_ net3 0.102f
C1979 _068_ a_6835_3968# 0.1f
C1980 VPWR ones[0] 0.288f
C1981 counter\[1\] _026_ 0.1f
C1982 _050_ _033_ 0.151f
C1983 _067_ clknet_1_0__leaf_clk 0.219f
C1984 counter\[1\] clknet_1_0__leaf_clk 0.261f
C1985 net9 _028_ 0.671f
C1986 VPWR _045_ 1.33f
C1987 a_6527_6263# net10 0.216f
C1988 _067_ _076_ 0.293f
C1989 _081_ _060_ 0.112f
C1990 net9 _035_ 0.133f
C1991 VPWR a_1589_5059# 0.207f
C1992 VPWR ones[2] 0.366f
C1993 VPWR _010_ 0.789f
C1994 _004_ a_8079_5162# 0.123f
C1995 VPWR _083_ 1.93f
C1996 _032_ _060_ 0.107f
C1997 _068_ _080_ 0.292f
C1998 net1 _022_ 0.23f
C1999 VPWR a_1846_2767# 0.282f
C2000 a_1547_10004# _007_ 0.129f
C2001 net7 _093_ 0.188f
C2002 _057_ _055_ 0.686f
C2003 net7 a_2603_9839# 0.251f
C2004 _005_ net2 1.76f
C2005 VPWR _043_ 2.79f
C2006 _012_ _083_ 2f
C2007 ones[8] ones[7] 0.124f
C2008 _036_ _045_ 0.75f
C2009 _056_ _028_ 0.177f
C2010 VPWR a_9551_5652# 0.25f
C2011 a_4234_9417# _029_ 0.171f
C2012 a_1407_10927# pulse 0.236f
C2013 _014_ net5 0.134f
C2014 counter\[10\] _084_ 0.476f
C2015 VPWR _004_ 0.653f
C2016 net13 _051_ 0.236f
C2017 _068_ counter\[0\] 0.336f
C2018 net9 net14 0.402f
C2019 _028_ _029_ 0.793f
C2020 _058_ net4 0.128f
C2021 a_4234_9417# _011_ 0.212f
C2022 _010_ a_3179_6031# 0.101f
C2023 _083_ net10 0.177f
C2024 _068_ counter\[8\] 0.181f
C2025 counter\[1\] counter\[2\] 2.32f
C2026 VPWR _074_ 1.32f
C2027 _070_ _074_ 0.129f
C2028 a_6007_8751# clknet_1_1__leaf_clk 0.301f
C2029 a_4035_7637# a_3939_7815# 0.311f
C2030 clk _046_ 0.151f
C2031 _059_ a_1589_5059# 0.203f
C2032 net7 a_9279_8725# 0.243f
C2033 _057_ net6 0.915f
C2034 _068_ _033_ 0.16f
C2035 _012_ _074_ 0.254f
C2036 a_4705_2767# _022_ 0.133f
C2037 counter\[2\] counter\[3\] 0.496f
C2038 VPWR counter\[9\] 2.13f
C2039 a_4517_2773# net3 0.163f
C2040 _084_ _060_ 0.34f
C2041 _004_ net10 0.463f
C2042 a_4351_2773# _023_ 0.114f
C2043 _056_ net14 0.147f
C2044 net6 net5 4.02f
C2045 a_4035_7637# VPWR 0.181f
C2046 net12 _027_ 0.263f
C2047 counter\[5\] _034_ 0.141f
C2048 VPWR a_5326_7093# 0.182f
C2049 net13 _014_ 0.155f
C2050 a_8352_9527# _033_ 0.122f
C2051 _039_ _049_ 0.619f
C2052 _074_ net10 0.235f
C2053 a_9711_2767# net5 0.123f
C2054 _071_ _060_ 0.107f
C2055 _066_ _081_ 0.896f
C2056 a_8307_10927# VPWR 0.228f
C2057 a_1573_2773# a_2014_2741# 0.119f
C2058 counter\[9\] _036_ 0.152f
C2059 _062_ _043_ 0.714f
C2060 _082_ _044_ 0.42f
C2061 VPWR a_4227_5161# 0.423f
C2062 VPWR a_9482_10383# 0.242f
C2063 rst a_1407_7119# 0.229f
C2064 _053_ VPWR 1.18f
C2065 _019_ _061_ 0.199f
C2066 VPWR _063_ 0.371f
C2067 a_7815_5461# clknet_1_1__leaf_clk 0.27f
C2068 _086_ net5 0.949f
C2069 ones[0] VGND 1.44f
C2070 ones[1] VGND 0.859f
C2071 ones[2] VGND 0.692f
C2072 ones[3] VGND 0.723f
C2073 ones[4] VGND 0.631f
C2074 ones[5] VGND 0.636f
C2075 clk VGND 2.03f
C2076 rst VGND 0.781f
C2077 ones[6] VGND 0.614f
C2078 ones[7] VGND 0.619f
C2079 ones[8] VGND 0.507f
C2080 ones[10] VGND 1.52f
C2081 ones[9] VGND 0.868f
C2082 ready VGND 1.93f
C2083 pulse VGND 1.06f
C2084 VPWR VGND 0.32p
C2085 a_10239_2223# VGND 0.229f
C2086 a_9963_2223# VGND 0.257f
C2087 a_5177_2487# VGND 0.244f
C2088 a_5077_2269# VGND 0.208f
C2089 a_1925_2473# VGND 0.329f
C2090 a_10075_3087# VGND 0.196f
C2091 a_9885_3087# VGND 0.165f
C2092 _088_ VGND 0.532f
C2093 a_7883_2767# VGND 0.294f
C2094 a_8051_2741# VGND 0.404f
C2095 a_7458_2767# VGND 0.245f
C2096 a_7626_2741# VGND 0.306f
C2097 a_7185_2773# VGND 0.456f
C2098 a_7019_2773# VGND 0.552f
C2099 a_6375_2775# VGND 0.381f
C2100 a_5215_2767# VGND 0.274f
C2101 a_5383_2741# VGND 0.47f
C2102 a_4790_2767# VGND 0.2f
C2103 a_4958_2741# VGND 0.248f
C2104 a_4517_2773# VGND 0.326f
C2105 a_4351_2773# VGND 0.476f
C2106 a_3932_2883# VGND 0.227f
C2107 a_2957_2999# VGND 0.239f
C2108 a_2271_2767# VGND 0.271f
C2109 a_2439_2741# VGND 0.38f
C2110 a_1846_2767# VGND 0.206f
C2111 a_2014_2741# VGND 0.248f
C2112 a_1573_2773# VGND 0.323f
C2113 a_1407_2773# VGND 0.515f
C2114 _024_ VGND 0.4f
C2115 a_5163_3311# VGND 0.241f
C2116 a_4719_3311# VGND 0.278f
C2117 a_10239_3311# VGND 0.268f
C2118 a_9544_3561# VGND 0.239f
C2119 a_7431_3285# VGND 0.242f
C2120 a_7255_3285# VGND 0.218f
C2121 a_6503_3677# VGND 0.26f
C2122 a_6671_3579# VGND 0.35f
C2123 a_6078_3677# VGND 0.205f
C2124 a_6246_3423# VGND 0.255f
C2125 a_5805_3311# VGND 0.335f
C2126 a_5639_3311# VGND 0.488f
C2127 _015_ VGND 2.54f
C2128 a_2971_3311# VGND 0.288f
C2129 a_7527_4087# VGND 0.298f
C2130 a_6835_3968# VGND 0.25f
C2131 a_4864_3829# VGND 0.365f
C2132 a_2419_4221# VGND 0.289f
C2133 a_1632_3971# VGND 0.215f
C2134 a_10239_4399# VGND 0.248f
C2135 a_7515_4765# VGND 0.282f
C2136 a_7683_4667# VGND 0.385f
C2137 a_7090_4765# VGND 0.199f
C2138 a_7258_4511# VGND 0.242f
C2139 a_6817_4399# VGND 0.306f
C2140 _017_ VGND 0.952f
C2141 a_6651_4399# VGND 0.474f
C2142 _077_ VGND 2.15f
C2143 a_2603_4405# VGND 0.331f
C2144 a_6375_4399# VGND 0.202f
C2145 a_6099_4399# VGND 0.244f
C2146 a_4903_4399# VGND 0.276f
C2147 a_3215_4551# VGND 0.268f
C2148 a_2795_4649# VGND 0.257f
C2149 _030_ VGND 0.56f
C2150 a_10011_5175# VGND 0.257f
C2151 a_8871_5321# VGND 0.256f
C2152 a_8942_5220# VGND 0.207f
C2153 a_8742_5065# VGND 0.33f
C2154 a_8735_5161# VGND 0.498f
C2155 a_8451_5175# VGND 0.275f
C2156 a_8355_5175# VGND 0.367f
C2157 a_8079_5162# VGND 0.211f
C2158 a_7123_5321# VGND 0.243f
C2159 a_7194_5220# VGND 0.2f
C2160 a_6994_5065# VGND 0.313f
C2161 a_6987_5161# VGND 0.472f
C2162 a_6703_5175# VGND 0.262f
C2163 a_6607_5175# VGND 0.36f
C2164 a_5779_5175# VGND 0.259f
C2165 a_4363_5321# VGND 0.252f
C2166 a_4434_5220# VGND 0.203f
C2167 a_4234_5065# VGND 0.31f
C2168 a_4227_5161# VGND 0.48f
C2169 a_3943_5175# VGND 0.266f
C2170 a_3847_5175# VGND 0.357f
C2171 a_2736_5059# VGND 0.25f
C2172 a_1589_5059# VGND 0.269f
C2173 _059_ VGND 3.22f
C2174 a_1489_4943# VGND 0.219f
C2175 _021_ VGND 0.315f
C2176 a_10239_5487# VGND 0.266f
C2177 a_9551_5652# VGND 0.244f
C2178 _052_ VGND 1.75f
C2179 _031_ VGND 2.49f
C2180 a_5316_5487# VGND 0.227f
C2181 _016_ VGND 0.479f
C2182 a_7951_5487# VGND 0.25f
C2183 a_8022_5461# VGND 0.198f
C2184 a_7815_5461# VGND 0.497f
C2185 a_7822_5761# VGND 0.316f
C2186 a_7531_5461# VGND 0.278f
C2187 a_7363_5461# VGND 0.444f
C2188 a_6546_5487# VGND 0.273f
C2189 _023_ VGND 2f
C2190 a_5915_5487# VGND 0.234f
C2191 a_5126_5487# VGND 0.249f
C2192 _038_ VGND 0.246f
C2193 a_4767_5652# VGND 0.225f
C2194 _001_ VGND 0.752f
C2195 a_2063_5487# VGND 0.266f
C2196 a_2134_5461# VGND 0.223f
C2197 a_1927_5461# VGND 0.544f
C2198 a_1934_5761# VGND 0.436f
C2199 a_1643_5461# VGND 0.274f
C2200 a_1475_5461# VGND 0.464f
C2201 _010_ VGND 0.581f
C2202 a_3368_6351# VGND 0.161f
C2203 a_3277_6351# VGND 0.125f
C2204 _067_ VGND 0.407f
C2205 a_9728_6147# VGND 0.234f
C2206 net8 VGND 2.13f
C2207 a_9275_6263# VGND 0.237f
C2208 a_8583_6397# VGND 0.238f
C2209 a_7975_6031# VGND 0.261f
C2210 a_8143_6005# VGND 0.338f
C2211 a_7550_6031# VGND 0.204f
C2212 a_7718_6005# VGND 0.247f
C2213 a_7277_6037# VGND 0.296f
C2214 _002_ VGND 0.405f
C2215 a_7111_6037# VGND 0.47f
C2216 a_6527_6263# VGND 0.229f
C2217 a_4053_6005# VGND 2.02f
C2218 a_3179_6031# VGND 0.204f
C2219 _090_ VGND 0.367f
C2220 a_2695_6144# VGND 0.267f
C2221 _065_ VGND 0.302f
C2222 a_1499_6031# VGND 0.238f
C2223 _032_ VGND 1.38f
C2224 _078_ VGND 1.21f
C2225 a_10239_6575# VGND 0.247f
C2226 net9 VGND 2.26f
C2227 _070_ VGND 1.42f
C2228 a_8263_6740# VGND 0.264f
C2229 a_5722_6575# VGND 2.06f
C2230 a_2051_6575# VGND 0.165f
C2231 counter\[10\] VGND 2.22f
C2232 _041_ VGND 0.647f
C2233 _083_ VGND 1.46f
C2234 _003_ VGND 2.33f
C2235 a_4363_6575# VGND 0.245f
C2236 a_4434_6549# VGND 0.204f
C2237 a_4227_6549# VGND 0.502f
C2238 a_4234_6849# VGND 0.317f
C2239 a_3943_6549# VGND 0.27f
C2240 a_3847_6727# VGND 0.353f
C2241 a_3247_6575# VGND 0.259f
C2242 a_2473_6549# VGND 0.287f
C2243 a_1669_6727# VGND 0.222f
C2244 a_10100_7351# VGND 0.204f
C2245 _091_ VGND 0.881f
C2246 a_9827_7351# VGND 0.235f
C2247 a_8022_7119# VGND 2.03f
C2248 clknet_0_clk VGND 2.27f
C2249 a_6375_7119# VGND 0.263f
C2250 a_5583_7119# VGND 0.259f
C2251 a_5751_7093# VGND 0.344f
C2252 a_5158_7119# VGND 0.221f
C2253 a_5326_7093# VGND 0.258f
C2254 a_4885_7125# VGND 0.301f
C2255 a_4719_7125# VGND 0.495f
C2256 _013_ VGND 0.399f
C2257 a_3259_7497# VGND 0.235f
C2258 a_3330_7396# VGND 0.192f
C2259 a_3130_7241# VGND 0.31f
C2260 a_3123_7337# VGND 0.494f
C2261 a_2839_7351# VGND 0.26f
C2262 a_2743_7351# VGND 0.377f
C2263 a_1407_7119# VGND 0.37f
C2264 _066_ VGND 1.78f
C2265 a_5684_7643# VGND 0.204f
C2266 a_10239_7663# VGND 0.262f
C2267 net10 VGND 2.82f
C2268 a_9306_7663# VGND 0.3f
C2269 _076_ VGND 0.64f
C2270 a_5411_7815# VGND 0.225f
C2271 _004_ VGND 0.875f
C2272 a_4455_7663# VGND 0.25f
C2273 a_4526_7637# VGND 0.205f
C2274 a_4319_7637# VGND 0.496f
C2275 a_4326_7937# VGND 0.337f
C2276 a_4035_7637# VGND 0.27f
C2277 a_3939_7815# VGND 0.373f
C2278 _064_ VGND 0.465f
C2279 _006_ VGND 0.476f
C2280 _048_ VGND 0.969f
C2281 _062_ VGND 0.79f
C2282 a_9919_8439# VGND 0.262f
C2283 _005_ VGND 2.77f
C2284 a_8963_8585# VGND 0.245f
C2285 a_9034_8484# VGND 0.194f
C2286 a_8834_8329# VGND 0.315f
C2287 a_8827_8425# VGND 0.47f
C2288 a_8543_8439# VGND 0.277f
C2289 a_8447_8439# VGND 0.376f
C2290 _079_ VGND 0.574f
C2291 a_5595_8426# VGND 0.26f
C2292 a_4627_8320# VGND 0.265f
C2293 _046_ VGND 0.471f
C2294 a_2271_8207# VGND 0.298f
C2295 a_2439_8181# VGND 0.516f
C2296 a_1846_8207# VGND 0.217f
C2297 a_2014_8181# VGND 0.257f
C2298 a_1573_8213# VGND 0.335f
C2299 _012_ VGND 2.56f
C2300 a_1407_8213# VGND 0.538f
C2301 _057_ VGND 1.35f
C2302 _058_ VGND 1.52f
C2303 _000_ VGND 0.573f
C2304 _009_ VGND 1.48f
C2305 a_9919_8903# VGND 0.249f
C2306 _037_ VGND 4f
C2307 a_9279_8725# VGND 0.258f
C2308 a_8215_8751# VGND 0.245f
C2309 _085_ VGND 1.34f
C2310 a_7895_8916# VGND 0.219f
C2311 _089_ VGND 2.85f
C2312 a_7619_8916# VGND 0.227f
C2313 a_6871_9117# VGND 0.251f
C2314 a_7039_9019# VGND 0.424f
C2315 a_6446_9117# VGND 0.202f
C2316 a_6614_8863# VGND 0.245f
C2317 a_6173_8751# VGND 0.296f
C2318 _014_ VGND 1.28f
C2319 a_6007_8751# VGND 0.484f
C2320 _075_ VGND 1.05f
C2321 _039_ VGND 2.74f
C2322 a_4338_8751# VGND 0.289f
C2323 counter\[5\] VGND 3.34f
C2324 a_2736_9001# VGND 0.259f
C2325 a_10239_9295# VGND 0.217f
C2326 a_9963_9295# VGND 0.223f
C2327 net2 VGND 5.66f
C2328 a_9088_9527# VGND 0.204f
C2329 _044_ VGND 0.512f
C2330 _033_ VGND 0.623f
C2331 a_8815_9527# VGND 0.239f
C2332 a_8352_9527# VGND 0.206f
C2333 _035_ VGND 0.923f
C2334 _036_ VGND 1.38f
C2335 _029_ VGND 0.469f
C2336 a_8079_9527# VGND 0.233f
C2337 _008_ VGND 0.305f
C2338 a_6939_9673# VGND 0.247f
C2339 a_7010_9572# VGND 0.203f
C2340 a_6810_9417# VGND 0.311f
C2341 a_6803_9513# VGND 0.493f
C2342 a_6519_9527# VGND 0.27f
C2343 a_6423_9527# VGND 0.354f
C2344 counter\[4\] VGND 2.72f
C2345 clknet_1_0__leaf_clk VGND 5.15f
C2346 a_4363_9673# VGND 0.238f
C2347 a_4434_9572# VGND 0.198f
C2348 a_4234_9417# VGND 0.357f
C2349 a_4227_9513# VGND 0.534f
C2350 a_3943_9527# VGND 0.271f
C2351 a_3775_9527# VGND 0.453f
C2352 a_3061_9411# VGND 0.249f
C2353 _027_ VGND 0.61f
C2354 a_2961_9295# VGND 0.202f
C2355 _022_ VGND 1.72f
C2356 a_2327_9295# VGND 0.259f
C2357 _045_ VGND 0.788f
C2358 a_1867_9295# VGND 0.263f
C2359 _054_ VGND 7.59f
C2360 _026_ VGND 3.64f
C2361 net11 VGND 3.57f
C2362 a_9655_9813# VGND 0.356f
C2363 a_7423_10205# VGND 0.282f
C2364 a_7591_10107# VGND 0.397f
C2365 a_6998_10205# VGND 0.195f
C2366 a_7166_9951# VGND 0.242f
C2367 a_6725_9839# VGND 0.325f
C2368 _018_ VGND 2.55f
C2369 a_6559_9839# VGND 0.479f
C2370 _081_ VGND 1.57f
C2371 _011_ VGND 0.536f
C2372 _050_ VGND 1.46f
C2373 _028_ VGND 4.14f
C2374 _049_ VGND 1.18f
C2375 _047_ VGND 0.855f
C2376 _055_ VGND 1.55f
C2377 _034_ VGND 0.843f
C2378 _007_ VGND 0.964f
C2379 a_6178_9839# VGND 0.286f
C2380 counter\[7\] VGND 3.87f
C2381 counter\[6\] VGND 2.36f
C2382 _074_ VGND 2.05f
C2383 _093_ VGND 2.03f
C2384 _092_ VGND 1.73f
C2385 a_4351_9839# VGND 0.244f
C2386 a_3970_9839# VGND 0.287f
C2387 _040_ VGND 1.6f
C2388 _042_ VGND 2.07f
C2389 a_3307_9991# VGND 0.261f
C2390 a_2603_9839# VGND 0.274f
C2391 net3 VGND 6.56f
C2392 net5 VGND 5.04f
C2393 net6 VGND 3.6f
C2394 net7 VGND 3.7f
C2395 _082_ VGND 1.85f
C2396 a_1547_10004# VGND 0.254f
C2397 _063_ VGND 1.09f
C2398 _053_ VGND 0.761f
C2399 _084_ VGND 0.975f
C2400 _073_ VGND 2.94f
C2401 _056_ VGND 1.6f
C2402 a_9907_10383# VGND 0.273f
C2403 a_10075_10357# VGND 0.368f
C2404 a_9482_10383# VGND 0.197f
C2405 a_9650_10357# VGND 0.256f
C2406 a_9209_10389# VGND 0.372f
C2407 _020_ VGND 0.44f
C2408 a_9043_10389# VGND 0.468f
C2409 a_8624_10499# VGND 0.218f
C2410 a_8307_10383# VGND 0.226f
C2411 a_7847_10383# VGND 0.218f
C2412 _051_ VGND 0.323f
C2413 a_7469_10703# VGND 0.239f
C2414 _025_ VGND 1.93f
C2415 net4 VGND 3.29f
C2416 _043_ VGND 2.22f
C2417 counter\[8\] VGND 3.61f
C2418 _080_ VGND 1.69f
C2419 _071_ VGND 0.667f
C2420 _072_ VGND 1.13f
C2421 a_2375_10615# VGND 0.281f
C2422 a_1665_10383# VGND 0.206f
C2423 a_1499_10383# VGND 0.283f
C2424 net12 VGND 6.67f
C2425 a_9815_11293# VGND 0.268f
C2426 a_9983_11195# VGND 0.45f
C2427 a_9390_11293# VGND 0.206f
C2428 a_9558_11039# VGND 0.245f
C2429 a_9117_10927# VGND 0.318f
C2430 _019_ VGND 1.84f
C2431 a_8951_10927# VGND 0.51f
C2432 clknet_1_1__leaf_clk VGND 4.53f
C2433 counter\[9\] VGND 1.86f
C2434 _086_ VGND 1.66f
C2435 _087_ VGND 1.63f
C2436 _068_ VGND 3.6f
C2437 _061_ VGND 0.756f
C2438 _069_ VGND 0.852f
C2439 net1 VGND 7.56f
C2440 a_8583_10927# VGND 0.215f
C2441 net13 VGND 3.19f
C2442 a_8307_10927# VGND 0.23f
C2443 net14 VGND 3.13f
C2444 a_5607_11079# VGND 0.267f
C2445 a_4043_10901# VGND 0.379f
C2446 a_3243_11293# VGND 0.226f
C2447 _060_ VGND 7.93f
C2448 a_3063_11293# VGND 0.231f
C2449 counter\[3\] VGND 1.42f
C2450 counter\[1\] VGND 6.38f
C2451 counter\[0\] VGND 4.01f
C2452 counter\[2\] VGND 3.76f
C2453 a_2472_10901# VGND 0.37f
C2454 a_1407_10927# VGND 0.387f
.ends

