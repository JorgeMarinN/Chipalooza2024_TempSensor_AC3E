magic
tech sky130A
magscale 1 2
timestamp 1712975979
<< checkpaint >>
rect -4008 -3980 4576 4524
<< poly >>
rect -76 199 118 265
<< locali >>
rect 218 215 416 265
<< viali >>
rect 462 219 496 253
<< metal1 >>
rect -76 496 644 592
rect 450 253 644 265
rect 450 219 462 253
rect 496 219 644 253
rect 450 199 644 219
rect -76 -48 644 48
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 54 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712864955
transform 1 0 330 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -38 0 1 0
box -38 -48 130 592
<< labels >>
rlabel poly -76 228 -76 228 7 VIN
port 1 w
rlabel metal1 644 234 644 234 3 VOUT
port 2 e
rlabel metal1 -76 -4 -76 -4 7 VSS
port 3 w
rlabel metal1 -76 540 -76 540 7 VDD
port 4 w
<< end >>
