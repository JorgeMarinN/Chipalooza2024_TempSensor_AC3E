magic
tech sky130A
magscale 1 2
timestamp 1713593032
<< error_s >>
rect -6001 19628 -5967 23948
rect 701 19628 735 23948
rect 1999 19628 2033 23948
rect 8701 19628 8735 23948
rect 9999 19628 10033 23948
rect 16701 19628 16735 23948
rect -6001 13856 -5967 18176
rect 701 13856 735 18176
rect 1999 13856 2033 18176
rect 8701 13856 8735 18176
rect 9999 13856 10033 18176
rect 16701 13856 16735 18176
rect -14853 9861 -14797 9881
rect -14773 9861 -14717 9881
rect -14885 9805 -14853 9861
rect -14797 9805 -14773 9861
rect -14717 9805 -14685 9861
rect -14853 9621 -14797 9805
rect -14773 9621 -14717 9805
rect -6001 8084 -5967 12404
rect 701 8084 735 12404
rect 1999 8084 2033 12404
rect 8701 8084 8735 12404
rect 9999 8084 10033 12404
rect 16701 8084 16735 12404
rect -6001 2312 -5967 6632
rect 701 2312 735 6632
rect 1999 2312 2033 6632
rect 8701 2312 8735 6632
rect 9999 2312 10033 6632
rect 16701 2312 16735 6632
rect -6001 -3460 -5967 860
rect 701 -3460 735 860
rect 1999 -3460 2033 860
rect 8701 -3460 8735 860
rect 9999 -3460 10033 860
rect 16701 -3460 16735 860
rect -8926 -14624 -8890 -14622
rect -8856 -14624 -8820 -14622
rect -7520 -14624 -7428 -14588
rect -6094 -14624 -6002 -14588
rect -4702 -14624 -4666 -14622
rect -4632 -14624 -4596 -14622
rect -8926 -14658 -7484 -14624
rect -7464 -14658 -6058 -14624
rect -6038 -14658 -4596 -14624
rect -8926 -17282 -8890 -14658
rect -8856 -17282 -8820 -14658
rect -7520 -14694 -7428 -14658
rect -6094 -14694 -6002 -14658
rect -7520 -17282 -7428 -17246
rect -6094 -17282 -6002 -17246
rect -4702 -17282 -4666 -14658
rect -4632 -17282 -4596 -14658
rect -8926 -17316 -7484 -17282
rect -7464 -17316 -6058 -17282
rect -6038 -17316 -4596 -17282
rect -8926 -17318 -8890 -17316
rect -8856 -17318 -8820 -17316
rect -7520 -17352 -7428 -17316
rect -6094 -17352 -6002 -17316
rect -4702 -17318 -4666 -17316
rect -4632 -17318 -4596 -17316
rect -14853 -18254 -14797 -18070
rect -14773 -18254 -14717 -18070
rect -14885 -18310 -14853 -18254
rect -14797 -18310 -14773 -18254
rect -14717 -18310 -14685 -18254
rect -14853 -18330 -14797 -18310
rect -14773 -18330 -14717 -18310
<< dnwell >>
rect -7630 10340 18381 24874
rect -30116 -18730 18381 10340
<< nwell >>
rect -7710 24668 18461 24954
rect -7710 10420 -7424 24668
rect -30196 10134 -7424 10420
rect -30196 -18524 -29910 10134
rect 18175 -18524 18461 24668
rect -30196 -18810 18461 -18524
<< nsubdiff >>
rect -6792 24858 -6622 24874
rect -6792 24818 -6762 24858
rect -6722 24818 -6688 24858
rect -6648 24818 -6622 24858
rect -6792 24784 -6622 24818
rect -6792 24744 -6762 24784
rect -6722 24744 -6688 24784
rect -6648 24744 -6622 24784
rect -6792 24714 -6622 24744
rect -4792 24858 -4622 24874
rect -4792 24818 -4762 24858
rect -4722 24818 -4688 24858
rect -4648 24818 -4622 24858
rect -4792 24784 -4622 24818
rect -4792 24744 -4762 24784
rect -4722 24744 -4688 24784
rect -4648 24744 -4622 24784
rect -4792 24714 -4622 24744
rect -2792 24858 -2622 24874
rect -2792 24818 -2762 24858
rect -2722 24818 -2688 24858
rect -2648 24818 -2622 24858
rect -2792 24784 -2622 24818
rect -2792 24744 -2762 24784
rect -2722 24744 -2688 24784
rect -2648 24744 -2622 24784
rect -2792 24714 -2622 24744
rect -792 24858 -622 24874
rect -792 24818 -762 24858
rect -722 24818 -688 24858
rect -648 24818 -622 24858
rect -792 24784 -622 24818
rect -792 24744 -762 24784
rect -722 24744 -688 24784
rect -648 24744 -622 24784
rect -792 24714 -622 24744
rect 1208 24858 1378 24874
rect 1208 24818 1238 24858
rect 1278 24818 1312 24858
rect 1352 24818 1378 24858
rect 1208 24784 1378 24818
rect 1208 24744 1238 24784
rect 1278 24744 1312 24784
rect 1352 24744 1378 24784
rect 1208 24714 1378 24744
rect 3208 24858 3378 24874
rect 3208 24818 3238 24858
rect 3278 24818 3312 24858
rect 3352 24818 3378 24858
rect 3208 24784 3378 24818
rect 3208 24744 3238 24784
rect 3278 24744 3312 24784
rect 3352 24744 3378 24784
rect 3208 24714 3378 24744
rect 5208 24858 5378 24874
rect 5208 24818 5238 24858
rect 5278 24818 5312 24858
rect 5352 24818 5378 24858
rect 5208 24784 5378 24818
rect 5208 24744 5238 24784
rect 5278 24744 5312 24784
rect 5352 24744 5378 24784
rect 5208 24714 5378 24744
rect 7208 24858 7378 24874
rect 7208 24818 7238 24858
rect 7278 24818 7312 24858
rect 7352 24818 7378 24858
rect 7208 24784 7378 24818
rect 7208 24744 7238 24784
rect 7278 24744 7312 24784
rect 7352 24744 7378 24784
rect 7208 24714 7378 24744
rect 9208 24858 9378 24874
rect 9208 24818 9238 24858
rect 9278 24818 9312 24858
rect 9352 24818 9378 24858
rect 9208 24784 9378 24818
rect 9208 24744 9238 24784
rect 9278 24744 9312 24784
rect 9352 24744 9378 24784
rect 9208 24714 9378 24744
rect 11208 24858 11378 24874
rect 11208 24818 11238 24858
rect 11278 24818 11312 24858
rect 11352 24818 11378 24858
rect 11208 24784 11378 24818
rect 11208 24744 11238 24784
rect 11278 24744 11312 24784
rect 11352 24744 11378 24784
rect 11208 24714 11378 24744
rect 13208 24858 13378 24874
rect 13208 24818 13238 24858
rect 13278 24818 13312 24858
rect 13352 24818 13378 24858
rect 13208 24784 13378 24818
rect 13208 24744 13238 24784
rect 13278 24744 13312 24784
rect 13352 24744 13378 24784
rect 13208 24714 13378 24744
rect 15208 24858 15378 24874
rect 15208 24818 15238 24858
rect 15278 24818 15312 24858
rect 15352 24818 15378 24858
rect 15208 24784 15378 24818
rect 15208 24744 15238 24784
rect 15278 24744 15312 24784
rect 15352 24744 15378 24784
rect 15208 24714 15378 24744
rect 17208 24858 17378 24874
rect 17208 24818 17238 24858
rect 17278 24818 17312 24858
rect 17352 24818 17378 24858
rect 17208 24784 17378 24818
rect 17208 24744 17238 24784
rect 17278 24744 17312 24784
rect 17352 24744 17378 24784
rect 17208 24714 17378 24744
rect -7630 24692 -7460 24708
rect -7630 24652 -7600 24692
rect -7560 24652 -7526 24692
rect -7486 24652 -7460 24692
rect -7630 24618 -7460 24652
rect -7630 24578 -7600 24618
rect -7560 24578 -7526 24618
rect -7486 24578 -7460 24618
rect -7630 24548 -7460 24578
rect 18212 23610 18380 23626
rect 18212 23570 18240 23610
rect 18280 23570 18314 23610
rect 18354 23570 18380 23610
rect 18212 23536 18380 23570
rect 18212 23496 18240 23536
rect 18280 23496 18314 23536
rect 18354 23496 18380 23536
rect 18212 23466 18380 23496
rect -7630 22692 -7460 22708
rect -7630 22652 -7600 22692
rect -7560 22652 -7526 22692
rect -7486 22652 -7460 22692
rect -7630 22618 -7460 22652
rect -7630 22578 -7600 22618
rect -7560 22578 -7526 22618
rect -7486 22578 -7460 22618
rect -7630 22548 -7460 22578
rect 18212 21610 18380 21626
rect 18212 21570 18240 21610
rect 18280 21570 18314 21610
rect 18354 21570 18380 21610
rect 18212 21536 18380 21570
rect 18212 21496 18240 21536
rect 18280 21496 18314 21536
rect 18354 21496 18380 21536
rect 18212 21466 18380 21496
rect -7630 20692 -7460 20708
rect -7630 20652 -7600 20692
rect -7560 20652 -7526 20692
rect -7486 20652 -7460 20692
rect -7630 20618 -7460 20652
rect -7630 20578 -7600 20618
rect -7560 20578 -7526 20618
rect -7486 20578 -7460 20618
rect -7630 20548 -7460 20578
rect 18212 19610 18380 19626
rect 18212 19570 18240 19610
rect 18280 19570 18314 19610
rect 18354 19570 18380 19610
rect 18212 19536 18380 19570
rect 18212 19496 18240 19536
rect 18280 19496 18314 19536
rect 18354 19496 18380 19536
rect 18212 19466 18380 19496
rect -7630 18692 -7460 18708
rect -7630 18652 -7600 18692
rect -7560 18652 -7526 18692
rect -7486 18652 -7460 18692
rect -7630 18618 -7460 18652
rect -7630 18578 -7600 18618
rect -7560 18578 -7526 18618
rect -7486 18578 -7460 18618
rect -7630 18548 -7460 18578
rect 18212 17610 18380 17626
rect 18212 17570 18240 17610
rect 18280 17570 18314 17610
rect 18354 17570 18380 17610
rect 18212 17536 18380 17570
rect 18212 17496 18240 17536
rect 18280 17496 18314 17536
rect 18354 17496 18380 17536
rect 18212 17466 18380 17496
rect -7630 16692 -7460 16708
rect -7630 16652 -7600 16692
rect -7560 16652 -7526 16692
rect -7486 16652 -7460 16692
rect -7630 16618 -7460 16652
rect -7630 16578 -7600 16618
rect -7560 16578 -7526 16618
rect -7486 16578 -7460 16618
rect -7630 16548 -7460 16578
rect 18212 15610 18380 15626
rect 18212 15570 18240 15610
rect 18280 15570 18314 15610
rect 18354 15570 18380 15610
rect 18212 15536 18380 15570
rect 18212 15496 18240 15536
rect 18280 15496 18314 15536
rect 18354 15496 18380 15536
rect 18212 15466 18380 15496
rect -7630 14692 -7460 14708
rect -7630 14652 -7600 14692
rect -7560 14652 -7526 14692
rect -7486 14652 -7460 14692
rect -7630 14618 -7460 14652
rect -7630 14578 -7600 14618
rect -7560 14578 -7526 14618
rect -7486 14578 -7460 14618
rect -7630 14548 -7460 14578
rect 18212 13610 18380 13626
rect 18212 13570 18240 13610
rect 18280 13570 18314 13610
rect 18354 13570 18380 13610
rect 18212 13536 18380 13570
rect 18212 13496 18240 13536
rect 18280 13496 18314 13536
rect 18354 13496 18380 13536
rect 18212 13466 18380 13496
rect -7630 12692 -7460 12708
rect -7630 12652 -7600 12692
rect -7560 12652 -7526 12692
rect -7486 12652 -7460 12692
rect -7630 12618 -7460 12652
rect -7630 12578 -7600 12618
rect -7560 12578 -7526 12618
rect -7486 12578 -7460 12618
rect -7630 12548 -7460 12578
rect 18212 11610 18380 11626
rect 18212 11570 18240 11610
rect 18280 11570 18314 11610
rect 18354 11570 18380 11610
rect 18212 11536 18380 11570
rect 18212 11496 18240 11536
rect 18280 11496 18314 11536
rect 18354 11496 18380 11536
rect 18212 11466 18380 11496
rect -7630 10692 -7460 10708
rect -7630 10652 -7600 10692
rect -7560 10652 -7526 10692
rect -7486 10652 -7460 10692
rect -7630 10618 -7460 10652
rect -7630 10578 -7600 10618
rect -7560 10578 -7526 10618
rect -7486 10578 -7460 10618
rect -7630 10548 -7460 10578
rect -29912 10324 -29742 10340
rect -29912 10284 -29882 10324
rect -29842 10284 -29808 10324
rect -29768 10284 -29742 10324
rect -29912 10250 -29742 10284
rect -29912 10210 -29882 10250
rect -29842 10210 -29808 10250
rect -29768 10210 -29742 10250
rect -29912 10180 -29742 10210
rect -27912 10324 -27742 10340
rect -27912 10284 -27882 10324
rect -27842 10284 -27808 10324
rect -27768 10284 -27742 10324
rect -27912 10250 -27742 10284
rect -27912 10210 -27882 10250
rect -27842 10210 -27808 10250
rect -27768 10210 -27742 10250
rect -27912 10180 -27742 10210
rect -25912 10324 -25742 10340
rect -25912 10284 -25882 10324
rect -25842 10284 -25808 10324
rect -25768 10284 -25742 10324
rect -25912 10250 -25742 10284
rect -25912 10210 -25882 10250
rect -25842 10210 -25808 10250
rect -25768 10210 -25742 10250
rect -25912 10180 -25742 10210
rect -23912 10324 -23742 10340
rect -23912 10284 -23882 10324
rect -23842 10284 -23808 10324
rect -23768 10284 -23742 10324
rect -23912 10250 -23742 10284
rect -23912 10210 -23882 10250
rect -23842 10210 -23808 10250
rect -23768 10210 -23742 10250
rect -23912 10180 -23742 10210
rect -21912 10324 -21742 10340
rect -21912 10284 -21882 10324
rect -21842 10284 -21808 10324
rect -21768 10284 -21742 10324
rect -21912 10250 -21742 10284
rect -21912 10210 -21882 10250
rect -21842 10210 -21808 10250
rect -21768 10210 -21742 10250
rect -21912 10180 -21742 10210
rect -19912 10324 -19742 10340
rect -19912 10284 -19882 10324
rect -19842 10284 -19808 10324
rect -19768 10284 -19742 10324
rect -19912 10250 -19742 10284
rect -19912 10210 -19882 10250
rect -19842 10210 -19808 10250
rect -19768 10210 -19742 10250
rect -19912 10180 -19742 10210
rect -17912 10324 -17742 10340
rect -17912 10284 -17882 10324
rect -17842 10284 -17808 10324
rect -17768 10284 -17742 10324
rect -17912 10250 -17742 10284
rect -17912 10210 -17882 10250
rect -17842 10210 -17808 10250
rect -17768 10210 -17742 10250
rect -17912 10180 -17742 10210
rect -15912 10324 -15742 10340
rect -15912 10284 -15882 10324
rect -15842 10284 -15808 10324
rect -15768 10284 -15742 10324
rect -15912 10250 -15742 10284
rect -15912 10210 -15882 10250
rect -15842 10210 -15808 10250
rect -15768 10210 -15742 10250
rect -15912 10180 -15742 10210
rect -13912 10324 -13742 10340
rect -13912 10284 -13882 10324
rect -13842 10284 -13808 10324
rect -13768 10284 -13742 10324
rect -13912 10250 -13742 10284
rect -13912 10210 -13882 10250
rect -13842 10210 -13808 10250
rect -13768 10210 -13742 10250
rect -13912 10180 -13742 10210
rect -11912 10324 -11742 10340
rect -11912 10284 -11882 10324
rect -11842 10284 -11808 10324
rect -11768 10284 -11742 10324
rect -11912 10250 -11742 10284
rect -11912 10210 -11882 10250
rect -11842 10210 -11808 10250
rect -11768 10210 -11742 10250
rect -11912 10180 -11742 10210
rect -9912 10324 -9742 10340
rect -9912 10284 -9882 10324
rect -9842 10284 -9808 10324
rect -9768 10284 -9742 10324
rect -9912 10250 -9742 10284
rect -9912 10210 -9882 10250
rect -9842 10210 -9808 10250
rect -9768 10210 -9742 10250
rect -9912 10180 -9742 10210
rect -7912 10324 -7742 10340
rect -7912 10284 -7882 10324
rect -7842 10284 -7808 10324
rect -7768 10284 -7742 10324
rect -7912 10250 -7742 10284
rect -7912 10210 -7882 10250
rect -7842 10210 -7808 10250
rect -7768 10210 -7742 10250
rect -7912 10180 -7742 10210
rect -30116 9622 -29946 9638
rect -30116 9582 -30086 9622
rect -30046 9582 -30012 9622
rect -29972 9582 -29946 9622
rect -30116 9548 -29946 9582
rect -30116 9508 -30086 9548
rect -30046 9508 -30012 9548
rect -29972 9508 -29946 9548
rect -30116 9478 -29946 9508
rect 18212 9610 18380 9626
rect 18212 9570 18240 9610
rect 18280 9570 18314 9610
rect 18354 9570 18380 9610
rect 18212 9536 18380 9570
rect 18212 9496 18240 9536
rect 18280 9496 18314 9536
rect 18354 9496 18380 9536
rect 18212 9466 18380 9496
rect -30116 7622 -29946 7638
rect -30116 7582 -30086 7622
rect -30046 7582 -30012 7622
rect -29972 7582 -29946 7622
rect -30116 7548 -29946 7582
rect -30116 7508 -30086 7548
rect -30046 7508 -30012 7548
rect -29972 7508 -29946 7548
rect -30116 7478 -29946 7508
rect 18212 7610 18380 7626
rect 18212 7570 18240 7610
rect 18280 7570 18314 7610
rect 18354 7570 18380 7610
rect 18212 7536 18380 7570
rect 18212 7496 18240 7536
rect 18280 7496 18314 7536
rect 18354 7496 18380 7536
rect 18212 7466 18380 7496
rect -30116 5622 -29946 5638
rect -30116 5582 -30086 5622
rect -30046 5582 -30012 5622
rect -29972 5582 -29946 5622
rect -30116 5548 -29946 5582
rect -30116 5508 -30086 5548
rect -30046 5508 -30012 5548
rect -29972 5508 -29946 5548
rect -30116 5478 -29946 5508
rect 18212 5610 18380 5626
rect 18212 5570 18240 5610
rect 18280 5570 18314 5610
rect 18354 5570 18380 5610
rect 18212 5536 18380 5570
rect 18212 5496 18240 5536
rect 18280 5496 18314 5536
rect 18354 5496 18380 5536
rect 18212 5466 18380 5496
rect -30116 3622 -29946 3638
rect -30116 3582 -30086 3622
rect -30046 3582 -30012 3622
rect -29972 3582 -29946 3622
rect -30116 3548 -29946 3582
rect -30116 3508 -30086 3548
rect -30046 3508 -30012 3548
rect -29972 3508 -29946 3548
rect -30116 3478 -29946 3508
rect 18212 3610 18380 3626
rect 18212 3570 18240 3610
rect 18280 3570 18314 3610
rect 18354 3570 18380 3610
rect 18212 3536 18380 3570
rect 18212 3496 18240 3536
rect 18280 3496 18314 3536
rect 18354 3496 18380 3536
rect 18212 3466 18380 3496
rect -30116 1622 -29946 1638
rect -30116 1582 -30086 1622
rect -30046 1582 -30012 1622
rect -29972 1582 -29946 1622
rect -30116 1548 -29946 1582
rect -30116 1508 -30086 1548
rect -30046 1508 -30012 1548
rect -29972 1508 -29946 1548
rect -30116 1478 -29946 1508
rect 18212 1610 18380 1626
rect 18212 1570 18240 1610
rect 18280 1570 18314 1610
rect 18354 1570 18380 1610
rect 18212 1536 18380 1570
rect 18212 1496 18240 1536
rect 18280 1496 18314 1536
rect 18354 1496 18380 1536
rect 18212 1466 18380 1496
rect -30116 -378 -29946 -362
rect -30116 -418 -30086 -378
rect -30046 -418 -30012 -378
rect -29972 -418 -29946 -378
rect -30116 -452 -29946 -418
rect -30116 -492 -30086 -452
rect -30046 -492 -30012 -452
rect -29972 -492 -29946 -452
rect -30116 -522 -29946 -492
rect 18212 -390 18380 -374
rect 18212 -430 18240 -390
rect 18280 -430 18314 -390
rect 18354 -430 18380 -390
rect 18212 -464 18380 -430
rect 18212 -504 18240 -464
rect 18280 -504 18314 -464
rect 18354 -504 18380 -464
rect 18212 -534 18380 -504
rect -30116 -2378 -29946 -2362
rect -30116 -2418 -30086 -2378
rect -30046 -2418 -30012 -2378
rect -29972 -2418 -29946 -2378
rect -30116 -2452 -29946 -2418
rect -30116 -2492 -30086 -2452
rect -30046 -2492 -30012 -2452
rect -29972 -2492 -29946 -2452
rect -30116 -2522 -29946 -2492
rect 18212 -2390 18380 -2374
rect 18212 -2430 18240 -2390
rect 18280 -2430 18314 -2390
rect 18354 -2430 18380 -2390
rect 18212 -2464 18380 -2430
rect 18212 -2504 18240 -2464
rect 18280 -2504 18314 -2464
rect 18354 -2504 18380 -2464
rect 18212 -2534 18380 -2504
rect -30116 -4378 -29946 -4362
rect -30116 -4418 -30086 -4378
rect -30046 -4418 -30012 -4378
rect -29972 -4418 -29946 -4378
rect -30116 -4452 -29946 -4418
rect -30116 -4492 -30086 -4452
rect -30046 -4492 -30012 -4452
rect -29972 -4492 -29946 -4452
rect -30116 -4522 -29946 -4492
rect 18212 -4390 18380 -4374
rect 18212 -4430 18240 -4390
rect 18280 -4430 18314 -4390
rect 18354 -4430 18380 -4390
rect 18212 -4464 18380 -4430
rect 18212 -4504 18240 -4464
rect 18280 -4504 18314 -4464
rect 18354 -4504 18380 -4464
rect 18212 -4534 18380 -4504
rect -30116 -6378 -29946 -6362
rect -30116 -6418 -30086 -6378
rect -30046 -6418 -30012 -6378
rect -29972 -6418 -29946 -6378
rect -30116 -6452 -29946 -6418
rect -30116 -6492 -30086 -6452
rect -30046 -6492 -30012 -6452
rect -29972 -6492 -29946 -6452
rect -30116 -6522 -29946 -6492
rect 18212 -6390 18380 -6374
rect 18212 -6430 18240 -6390
rect 18280 -6430 18314 -6390
rect 18354 -6430 18380 -6390
rect 18212 -6464 18380 -6430
rect 18212 -6504 18240 -6464
rect 18280 -6504 18314 -6464
rect 18354 -6504 18380 -6464
rect 18212 -6534 18380 -6504
rect -30116 -8378 -29946 -8362
rect -30116 -8418 -30086 -8378
rect -30046 -8418 -30012 -8378
rect -29972 -8418 -29946 -8378
rect -30116 -8452 -29946 -8418
rect -30116 -8492 -30086 -8452
rect -30046 -8492 -30012 -8452
rect -29972 -8492 -29946 -8452
rect -30116 -8522 -29946 -8492
rect 18212 -8390 18380 -8374
rect 18212 -8430 18240 -8390
rect 18280 -8430 18314 -8390
rect 18354 -8430 18380 -8390
rect 18212 -8464 18380 -8430
rect 18212 -8504 18240 -8464
rect 18280 -8504 18314 -8464
rect 18354 -8504 18380 -8464
rect 18212 -8534 18380 -8504
rect -30116 -10378 -29946 -10362
rect -30116 -10418 -30086 -10378
rect -30046 -10418 -30012 -10378
rect -29972 -10418 -29946 -10378
rect -30116 -10452 -29946 -10418
rect -30116 -10492 -30086 -10452
rect -30046 -10492 -30012 -10452
rect -29972 -10492 -29946 -10452
rect -30116 -10522 -29946 -10492
rect 18212 -10390 18380 -10374
rect 18212 -10430 18240 -10390
rect 18280 -10430 18314 -10390
rect 18354 -10430 18380 -10390
rect 18212 -10464 18380 -10430
rect 18212 -10504 18240 -10464
rect 18280 -10504 18314 -10464
rect 18354 -10504 18380 -10464
rect 18212 -10534 18380 -10504
rect -30116 -12378 -29946 -12362
rect -30116 -12418 -30086 -12378
rect -30046 -12418 -30012 -12378
rect -29972 -12418 -29946 -12378
rect -30116 -12452 -29946 -12418
rect -30116 -12492 -30086 -12452
rect -30046 -12492 -30012 -12452
rect -29972 -12492 -29946 -12452
rect -30116 -12522 -29946 -12492
rect 18212 -12390 18380 -12374
rect 18212 -12430 18240 -12390
rect 18280 -12430 18314 -12390
rect 18354 -12430 18380 -12390
rect 18212 -12464 18380 -12430
rect 18212 -12504 18240 -12464
rect 18280 -12504 18314 -12464
rect 18354 -12504 18380 -12464
rect 18212 -12534 18380 -12504
rect -30116 -14378 -29946 -14362
rect -30116 -14418 -30086 -14378
rect -30046 -14418 -30012 -14378
rect -29972 -14418 -29946 -14378
rect -30116 -14452 -29946 -14418
rect -30116 -14492 -30086 -14452
rect -30046 -14492 -30012 -14452
rect -29972 -14492 -29946 -14452
rect -30116 -14522 -29946 -14492
rect 18212 -14390 18380 -14374
rect 18212 -14430 18240 -14390
rect 18280 -14430 18314 -14390
rect 18354 -14430 18380 -14390
rect 18212 -14464 18380 -14430
rect 18212 -14504 18240 -14464
rect 18280 -14504 18314 -14464
rect 18354 -14504 18380 -14464
rect 18212 -14534 18380 -14504
rect -30116 -16378 -29946 -16362
rect -30116 -16418 -30086 -16378
rect -30046 -16418 -30012 -16378
rect -29972 -16418 -29946 -16378
rect -30116 -16452 -29946 -16418
rect -30116 -16492 -30086 -16452
rect -30046 -16492 -30012 -16452
rect -29972 -16492 -29946 -16452
rect -30116 -16522 -29946 -16492
rect 18212 -16390 18380 -16374
rect 18212 -16430 18240 -16390
rect 18280 -16430 18314 -16390
rect 18354 -16430 18380 -16390
rect 18212 -16464 18380 -16430
rect 18212 -16504 18240 -16464
rect 18280 -16504 18314 -16464
rect 18354 -16504 18380 -16464
rect 18212 -16534 18380 -16504
rect -30116 -18378 -29946 -18362
rect -30116 -18418 -30086 -18378
rect -30046 -18418 -30012 -18378
rect -29972 -18418 -29946 -18378
rect -30116 -18452 -29946 -18418
rect -30116 -18492 -30086 -18452
rect -30046 -18492 -30012 -18452
rect -29972 -18492 -29946 -18452
rect -30116 -18522 -29946 -18492
rect 18212 -18390 18380 -18374
rect 18212 -18430 18240 -18390
rect 18280 -18430 18314 -18390
rect 18354 -18430 18380 -18390
rect 18212 -18464 18380 -18430
rect 18212 -18504 18240 -18464
rect 18280 -18504 18314 -18464
rect 18354 -18504 18380 -18464
rect 18212 -18534 18380 -18504
rect -28942 -18582 -28774 -18566
rect -28942 -18622 -28914 -18582
rect -28874 -18622 -28840 -18582
rect -28800 -18622 -28774 -18582
rect -28942 -18656 -28774 -18622
rect -28942 -18696 -28914 -18656
rect -28874 -18696 -28840 -18656
rect -28800 -18696 -28774 -18656
rect -28942 -18726 -28774 -18696
rect -26942 -18582 -26774 -18566
rect -26942 -18622 -26914 -18582
rect -26874 -18622 -26840 -18582
rect -26800 -18622 -26774 -18582
rect -26942 -18656 -26774 -18622
rect -26942 -18696 -26914 -18656
rect -26874 -18696 -26840 -18656
rect -26800 -18696 -26774 -18656
rect -26942 -18726 -26774 -18696
rect -24942 -18582 -24774 -18566
rect -24942 -18622 -24914 -18582
rect -24874 -18622 -24840 -18582
rect -24800 -18622 -24774 -18582
rect -24942 -18656 -24774 -18622
rect -24942 -18696 -24914 -18656
rect -24874 -18696 -24840 -18656
rect -24800 -18696 -24774 -18656
rect -24942 -18726 -24774 -18696
rect -22942 -18582 -22774 -18566
rect -22942 -18622 -22914 -18582
rect -22874 -18622 -22840 -18582
rect -22800 -18622 -22774 -18582
rect -22942 -18656 -22774 -18622
rect -22942 -18696 -22914 -18656
rect -22874 -18696 -22840 -18656
rect -22800 -18696 -22774 -18656
rect -22942 -18726 -22774 -18696
rect -20942 -18582 -20774 -18566
rect -20942 -18622 -20914 -18582
rect -20874 -18622 -20840 -18582
rect -20800 -18622 -20774 -18582
rect -20942 -18656 -20774 -18622
rect -20942 -18696 -20914 -18656
rect -20874 -18696 -20840 -18656
rect -20800 -18696 -20774 -18656
rect -20942 -18726 -20774 -18696
rect -18942 -18582 -18774 -18566
rect -18942 -18622 -18914 -18582
rect -18874 -18622 -18840 -18582
rect -18800 -18622 -18774 -18582
rect -18942 -18656 -18774 -18622
rect -18942 -18696 -18914 -18656
rect -18874 -18696 -18840 -18656
rect -18800 -18696 -18774 -18656
rect -18942 -18726 -18774 -18696
rect -16942 -18582 -16774 -18566
rect -16942 -18622 -16914 -18582
rect -16874 -18622 -16840 -18582
rect -16800 -18622 -16774 -18582
rect -16942 -18656 -16774 -18622
rect -16942 -18696 -16914 -18656
rect -16874 -18696 -16840 -18656
rect -16800 -18696 -16774 -18656
rect -16942 -18726 -16774 -18696
rect -14942 -18582 -14774 -18566
rect -14942 -18622 -14914 -18582
rect -14874 -18622 -14840 -18582
rect -14800 -18622 -14774 -18582
rect -14942 -18656 -14774 -18622
rect -14942 -18696 -14914 -18656
rect -14874 -18696 -14840 -18656
rect -14800 -18696 -14774 -18656
rect -14942 -18726 -14774 -18696
rect -12942 -18582 -12774 -18566
rect -12942 -18622 -12914 -18582
rect -12874 -18622 -12840 -18582
rect -12800 -18622 -12774 -18582
rect -12942 -18656 -12774 -18622
rect -12942 -18696 -12914 -18656
rect -12874 -18696 -12840 -18656
rect -12800 -18696 -12774 -18656
rect -12942 -18726 -12774 -18696
rect -10942 -18582 -10774 -18566
rect -10942 -18622 -10914 -18582
rect -10874 -18622 -10840 -18582
rect -10800 -18622 -10774 -18582
rect -10942 -18656 -10774 -18622
rect -10942 -18696 -10914 -18656
rect -10874 -18696 -10840 -18656
rect -10800 -18696 -10774 -18656
rect -10942 -18726 -10774 -18696
rect -8942 -18582 -8774 -18566
rect -8942 -18622 -8914 -18582
rect -8874 -18622 -8840 -18582
rect -8800 -18622 -8774 -18582
rect -8942 -18656 -8774 -18622
rect -8942 -18696 -8914 -18656
rect -8874 -18696 -8840 -18656
rect -8800 -18696 -8774 -18656
rect -8942 -18726 -8774 -18696
rect -6942 -18582 -6774 -18566
rect -6942 -18622 -6914 -18582
rect -6874 -18622 -6840 -18582
rect -6800 -18622 -6774 -18582
rect -6942 -18656 -6774 -18622
rect -6942 -18696 -6914 -18656
rect -6874 -18696 -6840 -18656
rect -6800 -18696 -6774 -18656
rect -6942 -18726 -6774 -18696
rect -4942 -18582 -4774 -18566
rect -4942 -18622 -4914 -18582
rect -4874 -18622 -4840 -18582
rect -4800 -18622 -4774 -18582
rect -4942 -18656 -4774 -18622
rect -4942 -18696 -4914 -18656
rect -4874 -18696 -4840 -18656
rect -4800 -18696 -4774 -18656
rect -4942 -18726 -4774 -18696
rect -2942 -18582 -2774 -18566
rect -2942 -18622 -2914 -18582
rect -2874 -18622 -2840 -18582
rect -2800 -18622 -2774 -18582
rect -2942 -18656 -2774 -18622
rect -2942 -18696 -2914 -18656
rect -2874 -18696 -2840 -18656
rect -2800 -18696 -2774 -18656
rect -2942 -18726 -2774 -18696
rect -942 -18582 -774 -18566
rect -942 -18622 -914 -18582
rect -874 -18622 -840 -18582
rect -800 -18622 -774 -18582
rect -942 -18656 -774 -18622
rect -942 -18696 -914 -18656
rect -874 -18696 -840 -18656
rect -800 -18696 -774 -18656
rect -942 -18726 -774 -18696
rect 1058 -18582 1226 -18566
rect 1058 -18622 1086 -18582
rect 1126 -18622 1160 -18582
rect 1200 -18622 1226 -18582
rect 1058 -18656 1226 -18622
rect 1058 -18696 1086 -18656
rect 1126 -18696 1160 -18656
rect 1200 -18696 1226 -18656
rect 1058 -18726 1226 -18696
rect 3058 -18582 3226 -18566
rect 3058 -18622 3086 -18582
rect 3126 -18622 3160 -18582
rect 3200 -18622 3226 -18582
rect 3058 -18656 3226 -18622
rect 3058 -18696 3086 -18656
rect 3126 -18696 3160 -18656
rect 3200 -18696 3226 -18656
rect 3058 -18726 3226 -18696
rect 5058 -18582 5226 -18566
rect 5058 -18622 5086 -18582
rect 5126 -18622 5160 -18582
rect 5200 -18622 5226 -18582
rect 5058 -18656 5226 -18622
rect 5058 -18696 5086 -18656
rect 5126 -18696 5160 -18656
rect 5200 -18696 5226 -18656
rect 5058 -18726 5226 -18696
rect 7058 -18582 7226 -18566
rect 7058 -18622 7086 -18582
rect 7126 -18622 7160 -18582
rect 7200 -18622 7226 -18582
rect 7058 -18656 7226 -18622
rect 7058 -18696 7086 -18656
rect 7126 -18696 7160 -18656
rect 7200 -18696 7226 -18656
rect 7058 -18726 7226 -18696
rect 9058 -18582 9226 -18566
rect 9058 -18622 9086 -18582
rect 9126 -18622 9160 -18582
rect 9200 -18622 9226 -18582
rect 9058 -18656 9226 -18622
rect 9058 -18696 9086 -18656
rect 9126 -18696 9160 -18656
rect 9200 -18696 9226 -18656
rect 9058 -18726 9226 -18696
rect 11058 -18582 11226 -18566
rect 11058 -18622 11086 -18582
rect 11126 -18622 11160 -18582
rect 11200 -18622 11226 -18582
rect 11058 -18656 11226 -18622
rect 11058 -18696 11086 -18656
rect 11126 -18696 11160 -18656
rect 11200 -18696 11226 -18656
rect 11058 -18726 11226 -18696
rect 13058 -18582 13226 -18566
rect 13058 -18622 13086 -18582
rect 13126 -18622 13160 -18582
rect 13200 -18622 13226 -18582
rect 13058 -18656 13226 -18622
rect 13058 -18696 13086 -18656
rect 13126 -18696 13160 -18656
rect 13200 -18696 13226 -18656
rect 13058 -18726 13226 -18696
rect 15058 -18582 15226 -18566
rect 15058 -18622 15086 -18582
rect 15126 -18622 15160 -18582
rect 15200 -18622 15226 -18582
rect 15058 -18656 15226 -18622
rect 15058 -18696 15086 -18656
rect 15126 -18696 15160 -18656
rect 15200 -18696 15226 -18656
rect 15058 -18726 15226 -18696
rect 17058 -18582 17226 -18566
rect 17058 -18622 17086 -18582
rect 17126 -18622 17160 -18582
rect 17200 -18622 17226 -18582
rect 17058 -18656 17226 -18622
rect 17058 -18696 17086 -18656
rect 17126 -18696 17160 -18656
rect 17200 -18696 17226 -18656
rect 17058 -18726 17226 -18696
<< nsubdiffcont >>
rect -6762 24818 -6722 24858
rect -6688 24818 -6648 24858
rect -6762 24744 -6722 24784
rect -6688 24744 -6648 24784
rect -4762 24818 -4722 24858
rect -4688 24818 -4648 24858
rect -4762 24744 -4722 24784
rect -4688 24744 -4648 24784
rect -2762 24818 -2722 24858
rect -2688 24818 -2648 24858
rect -2762 24744 -2722 24784
rect -2688 24744 -2648 24784
rect -762 24818 -722 24858
rect -688 24818 -648 24858
rect -762 24744 -722 24784
rect -688 24744 -648 24784
rect 1238 24818 1278 24858
rect 1312 24818 1352 24858
rect 1238 24744 1278 24784
rect 1312 24744 1352 24784
rect 3238 24818 3278 24858
rect 3312 24818 3352 24858
rect 3238 24744 3278 24784
rect 3312 24744 3352 24784
rect 5238 24818 5278 24858
rect 5312 24818 5352 24858
rect 5238 24744 5278 24784
rect 5312 24744 5352 24784
rect 7238 24818 7278 24858
rect 7312 24818 7352 24858
rect 7238 24744 7278 24784
rect 7312 24744 7352 24784
rect 9238 24818 9278 24858
rect 9312 24818 9352 24858
rect 9238 24744 9278 24784
rect 9312 24744 9352 24784
rect 11238 24818 11278 24858
rect 11312 24818 11352 24858
rect 11238 24744 11278 24784
rect 11312 24744 11352 24784
rect 13238 24818 13278 24858
rect 13312 24818 13352 24858
rect 13238 24744 13278 24784
rect 13312 24744 13352 24784
rect 15238 24818 15278 24858
rect 15312 24818 15352 24858
rect 15238 24744 15278 24784
rect 15312 24744 15352 24784
rect 17238 24818 17278 24858
rect 17312 24818 17352 24858
rect 17238 24744 17278 24784
rect 17312 24744 17352 24784
rect -7600 24652 -7560 24692
rect -7526 24652 -7486 24692
rect -7600 24578 -7560 24618
rect -7526 24578 -7486 24618
rect 18240 23570 18280 23610
rect 18314 23570 18354 23610
rect 18240 23496 18280 23536
rect 18314 23496 18354 23536
rect -7600 22652 -7560 22692
rect -7526 22652 -7486 22692
rect -7600 22578 -7560 22618
rect -7526 22578 -7486 22618
rect 18240 21570 18280 21610
rect 18314 21570 18354 21610
rect 18240 21496 18280 21536
rect 18314 21496 18354 21536
rect -7600 20652 -7560 20692
rect -7526 20652 -7486 20692
rect -7600 20578 -7560 20618
rect -7526 20578 -7486 20618
rect 18240 19570 18280 19610
rect 18314 19570 18354 19610
rect 18240 19496 18280 19536
rect 18314 19496 18354 19536
rect -7600 18652 -7560 18692
rect -7526 18652 -7486 18692
rect -7600 18578 -7560 18618
rect -7526 18578 -7486 18618
rect 18240 17570 18280 17610
rect 18314 17570 18354 17610
rect 18240 17496 18280 17536
rect 18314 17496 18354 17536
rect -7600 16652 -7560 16692
rect -7526 16652 -7486 16692
rect -7600 16578 -7560 16618
rect -7526 16578 -7486 16618
rect 18240 15570 18280 15610
rect 18314 15570 18354 15610
rect 18240 15496 18280 15536
rect 18314 15496 18354 15536
rect -7600 14652 -7560 14692
rect -7526 14652 -7486 14692
rect -7600 14578 -7560 14618
rect -7526 14578 -7486 14618
rect 18240 13570 18280 13610
rect 18314 13570 18354 13610
rect 18240 13496 18280 13536
rect 18314 13496 18354 13536
rect -7600 12652 -7560 12692
rect -7526 12652 -7486 12692
rect -7600 12578 -7560 12618
rect -7526 12578 -7486 12618
rect 18240 11570 18280 11610
rect 18314 11570 18354 11610
rect 18240 11496 18280 11536
rect 18314 11496 18354 11536
rect -7600 10652 -7560 10692
rect -7526 10652 -7486 10692
rect -7600 10578 -7560 10618
rect -7526 10578 -7486 10618
rect -29882 10284 -29842 10324
rect -29808 10284 -29768 10324
rect -29882 10210 -29842 10250
rect -29808 10210 -29768 10250
rect -27882 10284 -27842 10324
rect -27808 10284 -27768 10324
rect -27882 10210 -27842 10250
rect -27808 10210 -27768 10250
rect -25882 10284 -25842 10324
rect -25808 10284 -25768 10324
rect -25882 10210 -25842 10250
rect -25808 10210 -25768 10250
rect -23882 10284 -23842 10324
rect -23808 10284 -23768 10324
rect -23882 10210 -23842 10250
rect -23808 10210 -23768 10250
rect -21882 10284 -21842 10324
rect -21808 10284 -21768 10324
rect -21882 10210 -21842 10250
rect -21808 10210 -21768 10250
rect -19882 10284 -19842 10324
rect -19808 10284 -19768 10324
rect -19882 10210 -19842 10250
rect -19808 10210 -19768 10250
rect -17882 10284 -17842 10324
rect -17808 10284 -17768 10324
rect -17882 10210 -17842 10250
rect -17808 10210 -17768 10250
rect -15882 10284 -15842 10324
rect -15808 10284 -15768 10324
rect -15882 10210 -15842 10250
rect -15808 10210 -15768 10250
rect -13882 10284 -13842 10324
rect -13808 10284 -13768 10324
rect -13882 10210 -13842 10250
rect -13808 10210 -13768 10250
rect -11882 10284 -11842 10324
rect -11808 10284 -11768 10324
rect -11882 10210 -11842 10250
rect -11808 10210 -11768 10250
rect -9882 10284 -9842 10324
rect -9808 10284 -9768 10324
rect -9882 10210 -9842 10250
rect -9808 10210 -9768 10250
rect -7882 10284 -7842 10324
rect -7808 10284 -7768 10324
rect -7882 10210 -7842 10250
rect -7808 10210 -7768 10250
rect -30086 9582 -30046 9622
rect -30012 9582 -29972 9622
rect -30086 9508 -30046 9548
rect -30012 9508 -29972 9548
rect 18240 9570 18280 9610
rect 18314 9570 18354 9610
rect 18240 9496 18280 9536
rect 18314 9496 18354 9536
rect -30086 7582 -30046 7622
rect -30012 7582 -29972 7622
rect -30086 7508 -30046 7548
rect -30012 7508 -29972 7548
rect 18240 7570 18280 7610
rect 18314 7570 18354 7610
rect 18240 7496 18280 7536
rect 18314 7496 18354 7536
rect -30086 5582 -30046 5622
rect -30012 5582 -29972 5622
rect -30086 5508 -30046 5548
rect -30012 5508 -29972 5548
rect 18240 5570 18280 5610
rect 18314 5570 18354 5610
rect 18240 5496 18280 5536
rect 18314 5496 18354 5536
rect -30086 3582 -30046 3622
rect -30012 3582 -29972 3622
rect -30086 3508 -30046 3548
rect -30012 3508 -29972 3548
rect 18240 3570 18280 3610
rect 18314 3570 18354 3610
rect 18240 3496 18280 3536
rect 18314 3496 18354 3536
rect -30086 1582 -30046 1622
rect -30012 1582 -29972 1622
rect -30086 1508 -30046 1548
rect -30012 1508 -29972 1548
rect 18240 1570 18280 1610
rect 18314 1570 18354 1610
rect 18240 1496 18280 1536
rect 18314 1496 18354 1536
rect -30086 -418 -30046 -378
rect -30012 -418 -29972 -378
rect -30086 -492 -30046 -452
rect -30012 -492 -29972 -452
rect 18240 -430 18280 -390
rect 18314 -430 18354 -390
rect 18240 -504 18280 -464
rect 18314 -504 18354 -464
rect -30086 -2418 -30046 -2378
rect -30012 -2418 -29972 -2378
rect -30086 -2492 -30046 -2452
rect -30012 -2492 -29972 -2452
rect 18240 -2430 18280 -2390
rect 18314 -2430 18354 -2390
rect 18240 -2504 18280 -2464
rect 18314 -2504 18354 -2464
rect -30086 -4418 -30046 -4378
rect -30012 -4418 -29972 -4378
rect -30086 -4492 -30046 -4452
rect -30012 -4492 -29972 -4452
rect 18240 -4430 18280 -4390
rect 18314 -4430 18354 -4390
rect 18240 -4504 18280 -4464
rect 18314 -4504 18354 -4464
rect -30086 -6418 -30046 -6378
rect -30012 -6418 -29972 -6378
rect -30086 -6492 -30046 -6452
rect -30012 -6492 -29972 -6452
rect 18240 -6430 18280 -6390
rect 18314 -6430 18354 -6390
rect 18240 -6504 18280 -6464
rect 18314 -6504 18354 -6464
rect -30086 -8418 -30046 -8378
rect -30012 -8418 -29972 -8378
rect -30086 -8492 -30046 -8452
rect -30012 -8492 -29972 -8452
rect 18240 -8430 18280 -8390
rect 18314 -8430 18354 -8390
rect 18240 -8504 18280 -8464
rect 18314 -8504 18354 -8464
rect -30086 -10418 -30046 -10378
rect -30012 -10418 -29972 -10378
rect -30086 -10492 -30046 -10452
rect -30012 -10492 -29972 -10452
rect 18240 -10430 18280 -10390
rect 18314 -10430 18354 -10390
rect 18240 -10504 18280 -10464
rect 18314 -10504 18354 -10464
rect -30086 -12418 -30046 -12378
rect -30012 -12418 -29972 -12378
rect -30086 -12492 -30046 -12452
rect -30012 -12492 -29972 -12452
rect 18240 -12430 18280 -12390
rect 18314 -12430 18354 -12390
rect 18240 -12504 18280 -12464
rect 18314 -12504 18354 -12464
rect -30086 -14418 -30046 -14378
rect -30012 -14418 -29972 -14378
rect -30086 -14492 -30046 -14452
rect -30012 -14492 -29972 -14452
rect 18240 -14430 18280 -14390
rect 18314 -14430 18354 -14390
rect 18240 -14504 18280 -14464
rect 18314 -14504 18354 -14464
rect -30086 -16418 -30046 -16378
rect -30012 -16418 -29972 -16378
rect -30086 -16492 -30046 -16452
rect -30012 -16492 -29972 -16452
rect 18240 -16430 18280 -16390
rect 18314 -16430 18354 -16390
rect 18240 -16504 18280 -16464
rect 18314 -16504 18354 -16464
rect -30086 -18418 -30046 -18378
rect -30012 -18418 -29972 -18378
rect -30086 -18492 -30046 -18452
rect -30012 -18492 -29972 -18452
rect 18240 -18430 18280 -18390
rect 18314 -18430 18354 -18390
rect 18240 -18504 18280 -18464
rect 18314 -18504 18354 -18464
rect -28914 -18622 -28874 -18582
rect -28840 -18622 -28800 -18582
rect -28914 -18696 -28874 -18656
rect -28840 -18696 -28800 -18656
rect -26914 -18622 -26874 -18582
rect -26840 -18622 -26800 -18582
rect -26914 -18696 -26874 -18656
rect -26840 -18696 -26800 -18656
rect -24914 -18622 -24874 -18582
rect -24840 -18622 -24800 -18582
rect -24914 -18696 -24874 -18656
rect -24840 -18696 -24800 -18656
rect -22914 -18622 -22874 -18582
rect -22840 -18622 -22800 -18582
rect -22914 -18696 -22874 -18656
rect -22840 -18696 -22800 -18656
rect -20914 -18622 -20874 -18582
rect -20840 -18622 -20800 -18582
rect -20914 -18696 -20874 -18656
rect -20840 -18696 -20800 -18656
rect -18914 -18622 -18874 -18582
rect -18840 -18622 -18800 -18582
rect -18914 -18696 -18874 -18656
rect -18840 -18696 -18800 -18656
rect -16914 -18622 -16874 -18582
rect -16840 -18622 -16800 -18582
rect -16914 -18696 -16874 -18656
rect -16840 -18696 -16800 -18656
rect -14914 -18622 -14874 -18582
rect -14840 -18622 -14800 -18582
rect -14914 -18696 -14874 -18656
rect -14840 -18696 -14800 -18656
rect -12914 -18622 -12874 -18582
rect -12840 -18622 -12800 -18582
rect -12914 -18696 -12874 -18656
rect -12840 -18696 -12800 -18656
rect -10914 -18622 -10874 -18582
rect -10840 -18622 -10800 -18582
rect -10914 -18696 -10874 -18656
rect -10840 -18696 -10800 -18656
rect -8914 -18622 -8874 -18582
rect -8840 -18622 -8800 -18582
rect -8914 -18696 -8874 -18656
rect -8840 -18696 -8800 -18656
rect -6914 -18622 -6874 -18582
rect -6840 -18622 -6800 -18582
rect -6914 -18696 -6874 -18656
rect -6840 -18696 -6800 -18656
rect -4914 -18622 -4874 -18582
rect -4840 -18622 -4800 -18582
rect -4914 -18696 -4874 -18656
rect -4840 -18696 -4800 -18656
rect -2914 -18622 -2874 -18582
rect -2840 -18622 -2800 -18582
rect -2914 -18696 -2874 -18656
rect -2840 -18696 -2800 -18656
rect -914 -18622 -874 -18582
rect -840 -18622 -800 -18582
rect -914 -18696 -874 -18656
rect -840 -18696 -800 -18656
rect 1086 -18622 1126 -18582
rect 1160 -18622 1200 -18582
rect 1086 -18696 1126 -18656
rect 1160 -18696 1200 -18656
rect 3086 -18622 3126 -18582
rect 3160 -18622 3200 -18582
rect 3086 -18696 3126 -18656
rect 3160 -18696 3200 -18656
rect 5086 -18622 5126 -18582
rect 5160 -18622 5200 -18582
rect 5086 -18696 5126 -18656
rect 5160 -18696 5200 -18656
rect 7086 -18622 7126 -18582
rect 7160 -18622 7200 -18582
rect 7086 -18696 7126 -18656
rect 7160 -18696 7200 -18656
rect 9086 -18622 9126 -18582
rect 9160 -18622 9200 -18582
rect 9086 -18696 9126 -18656
rect 9160 -18696 9200 -18656
rect 11086 -18622 11126 -18582
rect 11160 -18622 11200 -18582
rect 11086 -18696 11126 -18656
rect 11160 -18696 11200 -18656
rect 13086 -18622 13126 -18582
rect 13160 -18622 13200 -18582
rect 13086 -18696 13126 -18656
rect 13160 -18696 13200 -18656
rect 15086 -18622 15126 -18582
rect 15160 -18622 15200 -18582
rect 15086 -18696 15126 -18656
rect 15160 -18696 15200 -18656
rect 17086 -18622 17126 -18582
rect 17160 -18622 17200 -18582
rect 17086 -18696 17126 -18656
rect 17160 -18696 17200 -18656
<< locali >>
rect -7630 24858 18381 24874
rect -7630 24818 -6762 24858
rect -6722 24818 -6688 24858
rect -6648 24818 -4762 24858
rect -4722 24818 -4688 24858
rect -4648 24818 -2762 24858
rect -2722 24818 -2688 24858
rect -2648 24818 -762 24858
rect -722 24818 -688 24858
rect -648 24818 1238 24858
rect 1278 24818 1312 24858
rect 1352 24818 3238 24858
rect 3278 24818 3312 24858
rect 3352 24818 5238 24858
rect 5278 24818 5312 24858
rect 5352 24818 7238 24858
rect 7278 24818 7312 24858
rect 7352 24818 9238 24858
rect 9278 24818 9312 24858
rect 9352 24818 11238 24858
rect 11278 24818 11312 24858
rect 11352 24818 13238 24858
rect 13278 24818 13312 24858
rect 13352 24818 15238 24858
rect 15278 24818 15312 24858
rect 15352 24818 17238 24858
rect 17278 24818 17312 24858
rect 17352 24818 18381 24858
rect -7630 24784 18381 24818
rect -7630 24744 -6762 24784
rect -6722 24744 -6688 24784
rect -6648 24744 -4762 24784
rect -4722 24744 -4688 24784
rect -4648 24744 -2762 24784
rect -2722 24744 -2688 24784
rect -2648 24744 -762 24784
rect -722 24744 -688 24784
rect -648 24744 1238 24784
rect 1278 24744 1312 24784
rect 1352 24744 3238 24784
rect 3278 24744 3312 24784
rect 3352 24744 5238 24784
rect 5278 24744 5312 24784
rect 5352 24744 7238 24784
rect 7278 24744 7312 24784
rect 7352 24744 9238 24784
rect 9278 24744 9312 24784
rect 9352 24744 11238 24784
rect 11278 24744 11312 24784
rect 11352 24744 13238 24784
rect 13278 24744 13312 24784
rect 13352 24744 15238 24784
rect 15278 24744 15312 24784
rect 15352 24744 17238 24784
rect 17278 24744 17312 24784
rect 17352 24744 18381 24784
rect -7630 24692 18381 24744
rect -7630 24652 -7600 24692
rect -7560 24652 -7526 24692
rect -7486 24668 18381 24692
rect -7486 24652 -7424 24668
rect -7630 24618 -7424 24652
rect -7630 24578 -7600 24618
rect -7560 24578 -7526 24618
rect -7486 24578 -7424 24618
rect -7630 22692 -7424 24578
rect -7630 22652 -7600 22692
rect -7560 22652 -7526 22692
rect -7486 22652 -7424 22692
rect -7630 22618 -7424 22652
rect -7630 22578 -7600 22618
rect -7560 22578 -7526 22618
rect -7486 22578 -7424 22618
rect -7630 20692 -7424 22578
rect -7630 20652 -7600 20692
rect -7560 20652 -7526 20692
rect -7486 20652 -7424 20692
rect -7630 20618 -7424 20652
rect -7630 20578 -7600 20618
rect -7560 20578 -7526 20618
rect -7486 20578 -7424 20618
rect -7630 18692 -7424 20578
rect -7630 18652 -7600 18692
rect -7560 18652 -7526 18692
rect -7486 18652 -7424 18692
rect -7630 18618 -7424 18652
rect -7630 18578 -7600 18618
rect -7560 18578 -7526 18618
rect -7486 18578 -7424 18618
rect -7630 16692 -7424 18578
rect -7630 16652 -7600 16692
rect -7560 16652 -7526 16692
rect -7486 16652 -7424 16692
rect -7630 16618 -7424 16652
rect -7630 16578 -7600 16618
rect -7560 16578 -7526 16618
rect -7486 16578 -7424 16618
rect -7630 14692 -7424 16578
rect -7630 14652 -7600 14692
rect -7560 14652 -7526 14692
rect -7486 14652 -7424 14692
rect -7630 14618 -7424 14652
rect -7630 14578 -7600 14618
rect -7560 14578 -7526 14618
rect -7486 14578 -7424 14618
rect -7630 12692 -7424 14578
rect -7630 12652 -7600 12692
rect -7560 12652 -7526 12692
rect -7486 12652 -7424 12692
rect -7630 12618 -7424 12652
rect -7630 12578 -7600 12618
rect -7560 12578 -7526 12618
rect -7486 12578 -7424 12618
rect -7630 10692 -7424 12578
rect -7630 10652 -7600 10692
rect -7560 10652 -7526 10692
rect -7486 10652 -7424 10692
rect -7630 10618 -7424 10652
rect -7630 10578 -7600 10618
rect -7560 10578 -7526 10618
rect -7486 10578 -7424 10618
rect -7630 10340 -7424 10578
rect -30116 10324 -7424 10340
rect -30116 10284 -29882 10324
rect -29842 10284 -29808 10324
rect -29768 10284 -27882 10324
rect -27842 10284 -27808 10324
rect -27768 10284 -25882 10324
rect -25842 10284 -25808 10324
rect -25768 10284 -23882 10324
rect -23842 10284 -23808 10324
rect -23768 10284 -21882 10324
rect -21842 10284 -21808 10324
rect -21768 10284 -19882 10324
rect -19842 10284 -19808 10324
rect -19768 10284 -17882 10324
rect -17842 10284 -17808 10324
rect -17768 10284 -15882 10324
rect -15842 10284 -15808 10324
rect -15768 10284 -13882 10324
rect -13842 10284 -13808 10324
rect -13768 10284 -11882 10324
rect -11842 10284 -11808 10324
rect -11768 10284 -9882 10324
rect -9842 10284 -9808 10324
rect -9768 10284 -7882 10324
rect -7842 10284 -7808 10324
rect -7768 10284 -7424 10324
rect -30116 10250 -7424 10284
rect -30116 10210 -29882 10250
rect -29842 10210 -29808 10250
rect -29768 10210 -27882 10250
rect -27842 10210 -27808 10250
rect -27768 10210 -25882 10250
rect -25842 10210 -25808 10250
rect -25768 10210 -23882 10250
rect -23842 10210 -23808 10250
rect -23768 10210 -21882 10250
rect -21842 10210 -21808 10250
rect -21768 10210 -19882 10250
rect -19842 10210 -19808 10250
rect -19768 10210 -17882 10250
rect -17842 10210 -17808 10250
rect -17768 10210 -15882 10250
rect -15842 10210 -15808 10250
rect -15768 10210 -13882 10250
rect -13842 10210 -13808 10250
rect -13768 10210 -11882 10250
rect -11842 10210 -11808 10250
rect -11768 10210 -9882 10250
rect -9842 10210 -9808 10250
rect -9768 10210 -7882 10250
rect -7842 10210 -7808 10250
rect -7768 10210 -7424 10250
rect -30116 10134 -7424 10210
rect 18175 23610 18381 24668
rect 18175 23570 18240 23610
rect 18280 23570 18314 23610
rect 18354 23570 18381 23610
rect 18175 23536 18381 23570
rect 18175 23496 18240 23536
rect 18280 23496 18314 23536
rect 18354 23496 18381 23536
rect 18175 21610 18381 23496
rect 18175 21570 18240 21610
rect 18280 21570 18314 21610
rect 18354 21570 18381 21610
rect 18175 21536 18381 21570
rect 18175 21496 18240 21536
rect 18280 21496 18314 21536
rect 18354 21496 18381 21536
rect 18175 19610 18381 21496
rect 18175 19570 18240 19610
rect 18280 19570 18314 19610
rect 18354 19570 18381 19610
rect 18175 19536 18381 19570
rect 18175 19496 18240 19536
rect 18280 19496 18314 19536
rect 18354 19496 18381 19536
rect 18175 17610 18381 19496
rect 18175 17570 18240 17610
rect 18280 17570 18314 17610
rect 18354 17570 18381 17610
rect 18175 17536 18381 17570
rect 18175 17496 18240 17536
rect 18280 17496 18314 17536
rect 18354 17496 18381 17536
rect 18175 15610 18381 17496
rect 18175 15570 18240 15610
rect 18280 15570 18314 15610
rect 18354 15570 18381 15610
rect 18175 15536 18381 15570
rect 18175 15496 18240 15536
rect 18280 15496 18314 15536
rect 18354 15496 18381 15536
rect 18175 13610 18381 15496
rect 18175 13570 18240 13610
rect 18280 13570 18314 13610
rect 18354 13570 18381 13610
rect 18175 13536 18381 13570
rect 18175 13496 18240 13536
rect 18280 13496 18314 13536
rect 18354 13496 18381 13536
rect 18175 11610 18381 13496
rect 18175 11570 18240 11610
rect 18280 11570 18314 11610
rect 18354 11570 18381 11610
rect 18175 11536 18381 11570
rect 18175 11496 18240 11536
rect 18280 11496 18314 11536
rect 18354 11496 18381 11536
rect -30116 9622 -29910 10134
rect -30116 9582 -30086 9622
rect -30046 9582 -30012 9622
rect -29972 9582 -29910 9622
rect -30116 9548 -29910 9582
rect -30116 9508 -30086 9548
rect -30046 9508 -30012 9548
rect -29972 9508 -29910 9548
rect -30116 7622 -29910 9508
rect -30116 7582 -30086 7622
rect -30046 7582 -30012 7622
rect -29972 7582 -29910 7622
rect -30116 7548 -29910 7582
rect -30116 7508 -30086 7548
rect -30046 7508 -30012 7548
rect -29972 7508 -29910 7548
rect -30116 5622 -29910 7508
rect -30116 5582 -30086 5622
rect -30046 5582 -30012 5622
rect -29972 5582 -29910 5622
rect -30116 5548 -29910 5582
rect -30116 5508 -30086 5548
rect -30046 5508 -30012 5548
rect -29972 5508 -29910 5548
rect -30116 3622 -29910 5508
rect -30116 3582 -30086 3622
rect -30046 3582 -30012 3622
rect -29972 3582 -29910 3622
rect -30116 3548 -29910 3582
rect -30116 3508 -30086 3548
rect -30046 3508 -30012 3548
rect -29972 3508 -29910 3548
rect -30116 1622 -29910 3508
rect -30116 1582 -30086 1622
rect -30046 1582 -30012 1622
rect -29972 1582 -29910 1622
rect -30116 1548 -29910 1582
rect -30116 1508 -30086 1548
rect -30046 1508 -30012 1548
rect -29972 1508 -29910 1548
rect -30116 -378 -29910 1508
rect -30116 -418 -30086 -378
rect -30046 -418 -30012 -378
rect -29972 -418 -29910 -378
rect -30116 -452 -29910 -418
rect -30116 -492 -30086 -452
rect -30046 -492 -30012 -452
rect -29972 -492 -29910 -452
rect -30116 -2378 -29910 -492
rect -30116 -2418 -30086 -2378
rect -30046 -2418 -30012 -2378
rect -29972 -2418 -29910 -2378
rect -30116 -2452 -29910 -2418
rect -30116 -2492 -30086 -2452
rect -30046 -2492 -30012 -2452
rect -29972 -2492 -29910 -2452
rect -30116 -4378 -29910 -2492
rect -30116 -4418 -30086 -4378
rect -30046 -4418 -30012 -4378
rect -29972 -4418 -29910 -4378
rect -30116 -4452 -29910 -4418
rect -30116 -4492 -30086 -4452
rect -30046 -4492 -30012 -4452
rect -29972 -4492 -29910 -4452
rect -30116 -6378 -29910 -4492
rect -30116 -6418 -30086 -6378
rect -30046 -6418 -30012 -6378
rect -29972 -6418 -29910 -6378
rect -30116 -6452 -29910 -6418
rect -30116 -6492 -30086 -6452
rect -30046 -6492 -30012 -6452
rect -29972 -6492 -29910 -6452
rect -30116 -8378 -29910 -6492
rect -30116 -8418 -30086 -8378
rect -30046 -8418 -30012 -8378
rect -29972 -8418 -29910 -8378
rect -30116 -8452 -29910 -8418
rect -30116 -8492 -30086 -8452
rect -30046 -8492 -30012 -8452
rect -29972 -8492 -29910 -8452
rect -30116 -10378 -29910 -8492
rect -30116 -10418 -30086 -10378
rect -30046 -10418 -30012 -10378
rect -29972 -10418 -29910 -10378
rect -30116 -10452 -29910 -10418
rect -30116 -10492 -30086 -10452
rect -30046 -10492 -30012 -10452
rect -29972 -10492 -29910 -10452
rect -30116 -12378 -29910 -10492
rect -30116 -12418 -30086 -12378
rect -30046 -12418 -30012 -12378
rect -29972 -12418 -29910 -12378
rect -30116 -12452 -29910 -12418
rect -30116 -12492 -30086 -12452
rect -30046 -12492 -30012 -12452
rect -29972 -12492 -29910 -12452
rect -30116 -14378 -29910 -12492
rect -30116 -14418 -30086 -14378
rect -30046 -14418 -30012 -14378
rect -29972 -14418 -29910 -14378
rect -30116 -14452 -29910 -14418
rect -30116 -14492 -30086 -14452
rect -30046 -14492 -30012 -14452
rect -29972 -14492 -29910 -14452
rect -30116 -16378 -29910 -14492
rect -30116 -16418 -30086 -16378
rect -30046 -16418 -30012 -16378
rect -29972 -16418 -29910 -16378
rect -30116 -16452 -29910 -16418
rect -30116 -16492 -30086 -16452
rect -30046 -16492 -30012 -16452
rect -29972 -16492 -29910 -16452
rect -30116 -18378 -29910 -16492
rect -30116 -18418 -30086 -18378
rect -30046 -18418 -30012 -18378
rect -29972 -18418 -29910 -18378
rect -30116 -18452 -29910 -18418
rect -30116 -18492 -30086 -18452
rect -30046 -18492 -30012 -18452
rect -29972 -18492 -29910 -18452
rect -30116 -18524 -29910 -18492
rect 18175 9610 18381 11496
rect 18175 9570 18240 9610
rect 18280 9570 18314 9610
rect 18354 9570 18381 9610
rect 18175 9536 18381 9570
rect 18175 9496 18240 9536
rect 18280 9496 18314 9536
rect 18354 9496 18381 9536
rect 18175 7610 18381 9496
rect 18175 7570 18240 7610
rect 18280 7570 18314 7610
rect 18354 7570 18381 7610
rect 18175 7536 18381 7570
rect 18175 7496 18240 7536
rect 18280 7496 18314 7536
rect 18354 7496 18381 7536
rect 18175 5610 18381 7496
rect 18175 5570 18240 5610
rect 18280 5570 18314 5610
rect 18354 5570 18381 5610
rect 18175 5536 18381 5570
rect 18175 5496 18240 5536
rect 18280 5496 18314 5536
rect 18354 5496 18381 5536
rect 18175 3610 18381 5496
rect 18175 3570 18240 3610
rect 18280 3570 18314 3610
rect 18354 3570 18381 3610
rect 18175 3536 18381 3570
rect 18175 3496 18240 3536
rect 18280 3496 18314 3536
rect 18354 3496 18381 3536
rect 18175 1610 18381 3496
rect 18175 1570 18240 1610
rect 18280 1570 18314 1610
rect 18354 1570 18381 1610
rect 18175 1536 18381 1570
rect 18175 1496 18240 1536
rect 18280 1496 18314 1536
rect 18354 1496 18381 1536
rect 18175 -390 18381 1496
rect 18175 -430 18240 -390
rect 18280 -430 18314 -390
rect 18354 -430 18381 -390
rect 18175 -464 18381 -430
rect 18175 -504 18240 -464
rect 18280 -504 18314 -464
rect 18354 -504 18381 -464
rect 18175 -2390 18381 -504
rect 18175 -2430 18240 -2390
rect 18280 -2430 18314 -2390
rect 18354 -2430 18381 -2390
rect 18175 -2464 18381 -2430
rect 18175 -2504 18240 -2464
rect 18280 -2504 18314 -2464
rect 18354 -2504 18381 -2464
rect 18175 -4390 18381 -2504
rect 18175 -4430 18240 -4390
rect 18280 -4430 18314 -4390
rect 18354 -4430 18381 -4390
rect 18175 -4464 18381 -4430
rect 18175 -4504 18240 -4464
rect 18280 -4504 18314 -4464
rect 18354 -4504 18381 -4464
rect 18175 -6390 18381 -4504
rect 18175 -6430 18240 -6390
rect 18280 -6430 18314 -6390
rect 18354 -6430 18381 -6390
rect 18175 -6464 18381 -6430
rect 18175 -6504 18240 -6464
rect 18280 -6504 18314 -6464
rect 18354 -6504 18381 -6464
rect 18175 -8390 18381 -6504
rect 18175 -8430 18240 -8390
rect 18280 -8430 18314 -8390
rect 18354 -8430 18381 -8390
rect 18175 -8464 18381 -8430
rect 18175 -8504 18240 -8464
rect 18280 -8504 18314 -8464
rect 18354 -8504 18381 -8464
rect 18175 -10390 18381 -8504
rect 18175 -10430 18240 -10390
rect 18280 -10430 18314 -10390
rect 18354 -10430 18381 -10390
rect 18175 -10464 18381 -10430
rect 18175 -10504 18240 -10464
rect 18280 -10504 18314 -10464
rect 18354 -10504 18381 -10464
rect 18175 -12390 18381 -10504
rect 18175 -12430 18240 -12390
rect 18280 -12430 18314 -12390
rect 18354 -12430 18381 -12390
rect 18175 -12464 18381 -12430
rect 18175 -12504 18240 -12464
rect 18280 -12504 18314 -12464
rect 18354 -12504 18381 -12464
rect 18175 -14390 18381 -12504
rect 18175 -14430 18240 -14390
rect 18280 -14430 18314 -14390
rect 18354 -14430 18381 -14390
rect 18175 -14464 18381 -14430
rect 18175 -14504 18240 -14464
rect 18280 -14504 18314 -14464
rect 18354 -14504 18381 -14464
rect 18175 -16390 18381 -14504
rect 18175 -16430 18240 -16390
rect 18280 -16430 18314 -16390
rect 18354 -16430 18381 -16390
rect 18175 -16464 18381 -16430
rect 18175 -16504 18240 -16464
rect 18280 -16504 18314 -16464
rect 18354 -16504 18381 -16464
rect 18175 -18390 18381 -16504
rect 18175 -18430 18240 -18390
rect 18280 -18430 18314 -18390
rect 18354 -18430 18381 -18390
rect 18175 -18464 18381 -18430
rect 18175 -18504 18240 -18464
rect 18280 -18504 18314 -18464
rect 18354 -18504 18381 -18464
rect 18175 -18524 18381 -18504
rect -30116 -18582 18381 -18524
rect -30116 -18622 -28914 -18582
rect -28874 -18622 -28840 -18582
rect -28800 -18622 -26914 -18582
rect -26874 -18622 -26840 -18582
rect -26800 -18622 -24914 -18582
rect -24874 -18622 -24840 -18582
rect -24800 -18622 -22914 -18582
rect -22874 -18622 -22840 -18582
rect -22800 -18622 -20914 -18582
rect -20874 -18622 -20840 -18582
rect -20800 -18622 -18914 -18582
rect -18874 -18622 -18840 -18582
rect -18800 -18622 -16914 -18582
rect -16874 -18622 -16840 -18582
rect -16800 -18622 -14914 -18582
rect -14874 -18622 -14840 -18582
rect -14800 -18622 -12914 -18582
rect -12874 -18622 -12840 -18582
rect -12800 -18622 -10914 -18582
rect -10874 -18622 -10840 -18582
rect -10800 -18622 -8914 -18582
rect -8874 -18622 -8840 -18582
rect -8800 -18622 -6914 -18582
rect -6874 -18622 -6840 -18582
rect -6800 -18622 -4914 -18582
rect -4874 -18622 -4840 -18582
rect -4800 -18622 -2914 -18582
rect -2874 -18622 -2840 -18582
rect -2800 -18622 -914 -18582
rect -874 -18622 -840 -18582
rect -800 -18622 1086 -18582
rect 1126 -18622 1160 -18582
rect 1200 -18622 3086 -18582
rect 3126 -18622 3160 -18582
rect 3200 -18622 5086 -18582
rect 5126 -18622 5160 -18582
rect 5200 -18622 7086 -18582
rect 7126 -18622 7160 -18582
rect 7200 -18622 9086 -18582
rect 9126 -18622 9160 -18582
rect 9200 -18622 11086 -18582
rect 11126 -18622 11160 -18582
rect 11200 -18622 13086 -18582
rect 13126 -18622 13160 -18582
rect 13200 -18622 15086 -18582
rect 15126 -18622 15160 -18582
rect 15200 -18622 17086 -18582
rect 17126 -18622 17160 -18582
rect 17200 -18622 18381 -18582
rect -30116 -18656 18381 -18622
rect -30116 -18696 -28914 -18656
rect -28874 -18696 -28840 -18656
rect -28800 -18696 -26914 -18656
rect -26874 -18696 -26840 -18656
rect -26800 -18696 -24914 -18656
rect -24874 -18696 -24840 -18656
rect -24800 -18696 -22914 -18656
rect -22874 -18696 -22840 -18656
rect -22800 -18696 -20914 -18656
rect -20874 -18696 -20840 -18656
rect -20800 -18696 -18914 -18656
rect -18874 -18696 -18840 -18656
rect -18800 -18696 -16914 -18656
rect -16874 -18696 -16840 -18656
rect -16800 -18696 -14914 -18656
rect -14874 -18696 -14840 -18656
rect -14800 -18696 -12914 -18656
rect -12874 -18696 -12840 -18656
rect -12800 -18696 -10914 -18656
rect -10874 -18696 -10840 -18656
rect -10800 -18696 -8914 -18656
rect -8874 -18696 -8840 -18656
rect -8800 -18696 -6914 -18656
rect -6874 -18696 -6840 -18656
rect -6800 -18696 -4914 -18656
rect -4874 -18696 -4840 -18656
rect -4800 -18696 -2914 -18656
rect -2874 -18696 -2840 -18656
rect -2800 -18696 -914 -18656
rect -874 -18696 -840 -18656
rect -800 -18696 1086 -18656
rect 1126 -18696 1160 -18656
rect 1200 -18696 3086 -18656
rect 3126 -18696 3160 -18656
rect 3200 -18696 5086 -18656
rect 5126 -18696 5160 -18656
rect 5200 -18696 7086 -18656
rect 7126 -18696 7160 -18656
rect 7200 -18696 9086 -18656
rect 9126 -18696 9160 -18656
rect 9200 -18696 11086 -18656
rect 11126 -18696 11160 -18656
rect 11200 -18696 13086 -18656
rect 13126 -18696 13160 -18656
rect 13200 -18696 15086 -18656
rect 15126 -18696 15160 -18656
rect 15200 -18696 17086 -18656
rect 17126 -18696 17160 -18656
rect 17200 -18696 18381 -18656
rect -30116 -18730 18381 -18696
<< metal1 >>
rect -7630 24668 18381 24874
rect -7630 10340 -7424 24668
rect -30116 10134 -7424 10340
rect -30116 -18524 -29910 10134
rect -3328 -16710 -2408 -16590
rect -3328 -18017 -3208 -16710
rect -9902 -18083 -3208 -18017
rect 18175 -18524 18381 24668
rect -30116 -18730 18381 -18524
<< metal2 >>
rect -11563 -7342 -11363 -4237
rect -11563 -7462 -2412 -7342
rect -3208 -16710 -2408 -16590
use ONES_COUNTER  ONES_COUNTER_0
timestamp 1713593032
transform 1 0 -3101 0 1 -18207
box 0 824 11908 12912
use SDC  SDC_0
timestamp 1713593032
transform 1 0 19 0 1 -21
box -29735 -18309 17962 24495
<< end >>
