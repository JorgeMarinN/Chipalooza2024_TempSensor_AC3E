magic
tech sky130A
magscale 1 2
timestamp 1713593032
<< dnwell >>
rect -2206 -3414 2206 3414
<< nwell >>
rect -2286 3208 2286 3494
rect -2286 -3208 -2000 3208
rect 2000 -3208 2286 3208
rect -2286 -3494 2286 -3208
<< pwell >>
rect -1986 3050 1986 3182
rect -1986 -3182 1986 -3050
<< rpw >>
rect -2000 -3050 2000 3050
<< psubdiff >>
rect -1960 3154 1960 3156
rect -1960 3052 -1921 3154
rect 1921 3052 1960 3154
rect -1960 3050 1960 3052
rect -1960 -3052 1960 -3050
rect -1960 -3154 -1921 -3052
rect 1921 -3154 1960 -3052
rect -1960 -3156 1960 -3154
<< nsubdiff >>
rect -2160 3334 -2057 3368
rect -2023 3334 -1989 3368
rect -1955 3334 -1921 3368
rect -1887 3334 -1853 3368
rect -1819 3334 -1785 3368
rect -1751 3334 -1717 3368
rect -1683 3334 -1649 3368
rect -1615 3334 -1581 3368
rect -1547 3334 -1513 3368
rect -1479 3334 -1445 3368
rect -1411 3334 -1377 3368
rect -1343 3334 -1309 3368
rect -1275 3334 -1241 3368
rect -1207 3334 -1173 3368
rect -1139 3334 -1105 3368
rect -1071 3334 -1037 3368
rect -1003 3334 -969 3368
rect -935 3334 -901 3368
rect -867 3334 -833 3368
rect -799 3334 -765 3368
rect -731 3334 -697 3368
rect -663 3334 -629 3368
rect -595 3334 -561 3368
rect -527 3334 -493 3368
rect -459 3334 -425 3368
rect -391 3334 -357 3368
rect -323 3334 -289 3368
rect -255 3334 -221 3368
rect -187 3334 -153 3368
rect -119 3334 -85 3368
rect -51 3334 -17 3368
rect 17 3334 51 3368
rect 85 3334 119 3368
rect 153 3334 187 3368
rect 221 3334 255 3368
rect 289 3334 323 3368
rect 357 3334 391 3368
rect 425 3334 459 3368
rect 493 3334 527 3368
rect 561 3334 595 3368
rect 629 3334 663 3368
rect 697 3334 731 3368
rect 765 3334 799 3368
rect 833 3334 867 3368
rect 901 3334 935 3368
rect 969 3334 1003 3368
rect 1037 3334 1071 3368
rect 1105 3334 1139 3368
rect 1173 3334 1207 3368
rect 1241 3334 1275 3368
rect 1309 3334 1343 3368
rect 1377 3334 1411 3368
rect 1445 3334 1479 3368
rect 1513 3334 1547 3368
rect 1581 3334 1615 3368
rect 1649 3334 1683 3368
rect 1717 3334 1751 3368
rect 1785 3334 1819 3368
rect 1853 3334 1887 3368
rect 1921 3334 1955 3368
rect 1989 3334 2023 3368
rect 2057 3334 2160 3368
rect -2160 3213 -2126 3334
rect -2160 3145 -2126 3179
rect 2126 3213 2160 3334
rect -2160 3077 -2126 3111
rect 2126 3145 2160 3179
rect 2126 3077 2160 3111
rect -2160 3009 -2126 3043
rect -2160 2941 -2126 2975
rect -2160 2873 -2126 2907
rect -2160 2805 -2126 2839
rect -2160 2737 -2126 2771
rect -2160 2669 -2126 2703
rect -2160 2601 -2126 2635
rect -2160 2533 -2126 2567
rect -2160 2465 -2126 2499
rect -2160 2397 -2126 2431
rect -2160 2329 -2126 2363
rect -2160 2261 -2126 2295
rect -2160 2193 -2126 2227
rect -2160 2125 -2126 2159
rect -2160 2057 -2126 2091
rect -2160 1989 -2126 2023
rect -2160 1921 -2126 1955
rect -2160 1853 -2126 1887
rect -2160 1785 -2126 1819
rect -2160 1717 -2126 1751
rect -2160 1649 -2126 1683
rect -2160 1581 -2126 1615
rect -2160 1513 -2126 1547
rect -2160 1445 -2126 1479
rect -2160 1377 -2126 1411
rect -2160 1309 -2126 1343
rect -2160 1241 -2126 1275
rect -2160 1173 -2126 1207
rect -2160 1105 -2126 1139
rect -2160 1037 -2126 1071
rect -2160 969 -2126 1003
rect -2160 901 -2126 935
rect -2160 833 -2126 867
rect -2160 765 -2126 799
rect -2160 697 -2126 731
rect -2160 629 -2126 663
rect -2160 561 -2126 595
rect -2160 493 -2126 527
rect -2160 425 -2126 459
rect -2160 357 -2126 391
rect -2160 289 -2126 323
rect -2160 221 -2126 255
rect -2160 153 -2126 187
rect -2160 85 -2126 119
rect -2160 17 -2126 51
rect -2160 -51 -2126 -17
rect -2160 -119 -2126 -85
rect -2160 -187 -2126 -153
rect -2160 -255 -2126 -221
rect -2160 -323 -2126 -289
rect -2160 -391 -2126 -357
rect -2160 -459 -2126 -425
rect -2160 -527 -2126 -493
rect -2160 -595 -2126 -561
rect -2160 -663 -2126 -629
rect -2160 -731 -2126 -697
rect -2160 -799 -2126 -765
rect -2160 -867 -2126 -833
rect -2160 -935 -2126 -901
rect -2160 -1003 -2126 -969
rect -2160 -1071 -2126 -1037
rect -2160 -1139 -2126 -1105
rect -2160 -1207 -2126 -1173
rect -2160 -1275 -2126 -1241
rect -2160 -1343 -2126 -1309
rect -2160 -1411 -2126 -1377
rect -2160 -1479 -2126 -1445
rect -2160 -1547 -2126 -1513
rect -2160 -1615 -2126 -1581
rect -2160 -1683 -2126 -1649
rect -2160 -1751 -2126 -1717
rect -2160 -1819 -2126 -1785
rect -2160 -1887 -2126 -1853
rect -2160 -1955 -2126 -1921
rect -2160 -2023 -2126 -1989
rect -2160 -2091 -2126 -2057
rect -2160 -2159 -2126 -2125
rect -2160 -2227 -2126 -2193
rect -2160 -2295 -2126 -2261
rect -2160 -2363 -2126 -2329
rect -2160 -2431 -2126 -2397
rect -2160 -2499 -2126 -2465
rect -2160 -2567 -2126 -2533
rect -2160 -2635 -2126 -2601
rect -2160 -2703 -2126 -2669
rect -2160 -2771 -2126 -2737
rect -2160 -2839 -2126 -2805
rect -2160 -2907 -2126 -2873
rect -2160 -2975 -2126 -2941
rect -2160 -3043 -2126 -3009
rect 2126 3009 2160 3043
rect 2126 2941 2160 2975
rect 2126 2873 2160 2907
rect 2126 2805 2160 2839
rect 2126 2737 2160 2771
rect 2126 2669 2160 2703
rect 2126 2601 2160 2635
rect 2126 2533 2160 2567
rect 2126 2465 2160 2499
rect 2126 2397 2160 2431
rect 2126 2329 2160 2363
rect 2126 2261 2160 2295
rect 2126 2193 2160 2227
rect 2126 2125 2160 2159
rect 2126 2057 2160 2091
rect 2126 1989 2160 2023
rect 2126 1921 2160 1955
rect 2126 1853 2160 1887
rect 2126 1785 2160 1819
rect 2126 1717 2160 1751
rect 2126 1649 2160 1683
rect 2126 1581 2160 1615
rect 2126 1513 2160 1547
rect 2126 1445 2160 1479
rect 2126 1377 2160 1411
rect 2126 1309 2160 1343
rect 2126 1241 2160 1275
rect 2126 1173 2160 1207
rect 2126 1105 2160 1139
rect 2126 1037 2160 1071
rect 2126 969 2160 1003
rect 2126 901 2160 935
rect 2126 833 2160 867
rect 2126 765 2160 799
rect 2126 697 2160 731
rect 2126 629 2160 663
rect 2126 561 2160 595
rect 2126 493 2160 527
rect 2126 425 2160 459
rect 2126 357 2160 391
rect 2126 289 2160 323
rect 2126 221 2160 255
rect 2126 153 2160 187
rect 2126 85 2160 119
rect 2126 17 2160 51
rect 2126 -51 2160 -17
rect 2126 -119 2160 -85
rect 2126 -187 2160 -153
rect 2126 -255 2160 -221
rect 2126 -323 2160 -289
rect 2126 -391 2160 -357
rect 2126 -459 2160 -425
rect 2126 -527 2160 -493
rect 2126 -595 2160 -561
rect 2126 -663 2160 -629
rect 2126 -731 2160 -697
rect 2126 -799 2160 -765
rect 2126 -867 2160 -833
rect 2126 -935 2160 -901
rect 2126 -1003 2160 -969
rect 2126 -1071 2160 -1037
rect 2126 -1139 2160 -1105
rect 2126 -1207 2160 -1173
rect 2126 -1275 2160 -1241
rect 2126 -1343 2160 -1309
rect 2126 -1411 2160 -1377
rect 2126 -1479 2160 -1445
rect 2126 -1547 2160 -1513
rect 2126 -1615 2160 -1581
rect 2126 -1683 2160 -1649
rect 2126 -1751 2160 -1717
rect 2126 -1819 2160 -1785
rect 2126 -1887 2160 -1853
rect 2126 -1955 2160 -1921
rect 2126 -2023 2160 -1989
rect 2126 -2091 2160 -2057
rect 2126 -2159 2160 -2125
rect 2126 -2227 2160 -2193
rect 2126 -2295 2160 -2261
rect 2126 -2363 2160 -2329
rect 2126 -2431 2160 -2397
rect 2126 -2499 2160 -2465
rect 2126 -2567 2160 -2533
rect 2126 -2635 2160 -2601
rect 2126 -2703 2160 -2669
rect 2126 -2771 2160 -2737
rect 2126 -2839 2160 -2805
rect 2126 -2907 2160 -2873
rect 2126 -2975 2160 -2941
rect 2126 -3043 2160 -3009
rect -2160 -3111 -2126 -3077
rect -2160 -3179 -2126 -3145
rect 2126 -3111 2160 -3077
rect -2160 -3334 -2126 -3213
rect 2126 -3179 2160 -3145
rect 2126 -3334 2160 -3213
rect -2160 -3368 -2057 -3334
rect -2023 -3368 -1989 -3334
rect -1955 -3368 -1921 -3334
rect -1887 -3368 -1853 -3334
rect -1819 -3368 -1785 -3334
rect -1751 -3368 -1717 -3334
rect -1683 -3368 -1649 -3334
rect -1615 -3368 -1581 -3334
rect -1547 -3368 -1513 -3334
rect -1479 -3368 -1445 -3334
rect -1411 -3368 -1377 -3334
rect -1343 -3368 -1309 -3334
rect -1275 -3368 -1241 -3334
rect -1207 -3368 -1173 -3334
rect -1139 -3368 -1105 -3334
rect -1071 -3368 -1037 -3334
rect -1003 -3368 -969 -3334
rect -935 -3368 -901 -3334
rect -867 -3368 -833 -3334
rect -799 -3368 -765 -3334
rect -731 -3368 -697 -3334
rect -663 -3368 -629 -3334
rect -595 -3368 -561 -3334
rect -527 -3368 -493 -3334
rect -459 -3368 -425 -3334
rect -391 -3368 -357 -3334
rect -323 -3368 -289 -3334
rect -255 -3368 -221 -3334
rect -187 -3368 -153 -3334
rect -119 -3368 -85 -3334
rect -51 -3368 -17 -3334
rect 17 -3368 51 -3334
rect 85 -3368 119 -3334
rect 153 -3368 187 -3334
rect 221 -3368 255 -3334
rect 289 -3368 323 -3334
rect 357 -3368 391 -3334
rect 425 -3368 459 -3334
rect 493 -3368 527 -3334
rect 561 -3368 595 -3334
rect 629 -3368 663 -3334
rect 697 -3368 731 -3334
rect 765 -3368 799 -3334
rect 833 -3368 867 -3334
rect 901 -3368 935 -3334
rect 969 -3368 1003 -3334
rect 1037 -3368 1071 -3334
rect 1105 -3368 1139 -3334
rect 1173 -3368 1207 -3334
rect 1241 -3368 1275 -3334
rect 1309 -3368 1343 -3334
rect 1377 -3368 1411 -3334
rect 1445 -3368 1479 -3334
rect 1513 -3368 1547 -3334
rect 1581 -3368 1615 -3334
rect 1649 -3368 1683 -3334
rect 1717 -3368 1751 -3334
rect 1785 -3368 1819 -3334
rect 1853 -3368 1887 -3334
rect 1921 -3368 1955 -3334
rect 1989 -3368 2023 -3334
rect 2057 -3368 2160 -3334
<< psubdiffcont >>
rect -1921 3052 1921 3154
rect -1921 -3154 1921 -3052
<< nsubdiffcont >>
rect -2057 3334 -2023 3368
rect -1989 3334 -1955 3368
rect -1921 3334 -1887 3368
rect -1853 3334 -1819 3368
rect -1785 3334 -1751 3368
rect -1717 3334 -1683 3368
rect -1649 3334 -1615 3368
rect -1581 3334 -1547 3368
rect -1513 3334 -1479 3368
rect -1445 3334 -1411 3368
rect -1377 3334 -1343 3368
rect -1309 3334 -1275 3368
rect -1241 3334 -1207 3368
rect -1173 3334 -1139 3368
rect -1105 3334 -1071 3368
rect -1037 3334 -1003 3368
rect -969 3334 -935 3368
rect -901 3334 -867 3368
rect -833 3334 -799 3368
rect -765 3334 -731 3368
rect -697 3334 -663 3368
rect -629 3334 -595 3368
rect -561 3334 -527 3368
rect -493 3334 -459 3368
rect -425 3334 -391 3368
rect -357 3334 -323 3368
rect -289 3334 -255 3368
rect -221 3334 -187 3368
rect -153 3334 -119 3368
rect -85 3334 -51 3368
rect -17 3334 17 3368
rect 51 3334 85 3368
rect 119 3334 153 3368
rect 187 3334 221 3368
rect 255 3334 289 3368
rect 323 3334 357 3368
rect 391 3334 425 3368
rect 459 3334 493 3368
rect 527 3334 561 3368
rect 595 3334 629 3368
rect 663 3334 697 3368
rect 731 3334 765 3368
rect 799 3334 833 3368
rect 867 3334 901 3368
rect 935 3334 969 3368
rect 1003 3334 1037 3368
rect 1071 3334 1105 3368
rect 1139 3334 1173 3368
rect 1207 3334 1241 3368
rect 1275 3334 1309 3368
rect 1343 3334 1377 3368
rect 1411 3334 1445 3368
rect 1479 3334 1513 3368
rect 1547 3334 1581 3368
rect 1615 3334 1649 3368
rect 1683 3334 1717 3368
rect 1751 3334 1785 3368
rect 1819 3334 1853 3368
rect 1887 3334 1921 3368
rect 1955 3334 1989 3368
rect 2023 3334 2057 3368
rect -2160 3179 -2126 3213
rect 2126 3179 2160 3213
rect -2160 3111 -2126 3145
rect -2160 3043 -2126 3077
rect 2126 3111 2160 3145
rect -2160 2975 -2126 3009
rect -2160 2907 -2126 2941
rect -2160 2839 -2126 2873
rect -2160 2771 -2126 2805
rect -2160 2703 -2126 2737
rect -2160 2635 -2126 2669
rect -2160 2567 -2126 2601
rect -2160 2499 -2126 2533
rect -2160 2431 -2126 2465
rect -2160 2363 -2126 2397
rect -2160 2295 -2126 2329
rect -2160 2227 -2126 2261
rect -2160 2159 -2126 2193
rect -2160 2091 -2126 2125
rect -2160 2023 -2126 2057
rect -2160 1955 -2126 1989
rect -2160 1887 -2126 1921
rect -2160 1819 -2126 1853
rect -2160 1751 -2126 1785
rect -2160 1683 -2126 1717
rect -2160 1615 -2126 1649
rect -2160 1547 -2126 1581
rect -2160 1479 -2126 1513
rect -2160 1411 -2126 1445
rect -2160 1343 -2126 1377
rect -2160 1275 -2126 1309
rect -2160 1207 -2126 1241
rect -2160 1139 -2126 1173
rect -2160 1071 -2126 1105
rect -2160 1003 -2126 1037
rect -2160 935 -2126 969
rect -2160 867 -2126 901
rect -2160 799 -2126 833
rect -2160 731 -2126 765
rect -2160 663 -2126 697
rect -2160 595 -2126 629
rect -2160 527 -2126 561
rect -2160 459 -2126 493
rect -2160 391 -2126 425
rect -2160 323 -2126 357
rect -2160 255 -2126 289
rect -2160 187 -2126 221
rect -2160 119 -2126 153
rect -2160 51 -2126 85
rect -2160 -17 -2126 17
rect -2160 -85 -2126 -51
rect -2160 -153 -2126 -119
rect -2160 -221 -2126 -187
rect -2160 -289 -2126 -255
rect -2160 -357 -2126 -323
rect -2160 -425 -2126 -391
rect -2160 -493 -2126 -459
rect -2160 -561 -2126 -527
rect -2160 -629 -2126 -595
rect -2160 -697 -2126 -663
rect -2160 -765 -2126 -731
rect -2160 -833 -2126 -799
rect -2160 -901 -2126 -867
rect -2160 -969 -2126 -935
rect -2160 -1037 -2126 -1003
rect -2160 -1105 -2126 -1071
rect -2160 -1173 -2126 -1139
rect -2160 -1241 -2126 -1207
rect -2160 -1309 -2126 -1275
rect -2160 -1377 -2126 -1343
rect -2160 -1445 -2126 -1411
rect -2160 -1513 -2126 -1479
rect -2160 -1581 -2126 -1547
rect -2160 -1649 -2126 -1615
rect -2160 -1717 -2126 -1683
rect -2160 -1785 -2126 -1751
rect -2160 -1853 -2126 -1819
rect -2160 -1921 -2126 -1887
rect -2160 -1989 -2126 -1955
rect -2160 -2057 -2126 -2023
rect -2160 -2125 -2126 -2091
rect -2160 -2193 -2126 -2159
rect -2160 -2261 -2126 -2227
rect -2160 -2329 -2126 -2295
rect -2160 -2397 -2126 -2363
rect -2160 -2465 -2126 -2431
rect -2160 -2533 -2126 -2499
rect -2160 -2601 -2126 -2567
rect -2160 -2669 -2126 -2635
rect -2160 -2737 -2126 -2703
rect -2160 -2805 -2126 -2771
rect -2160 -2873 -2126 -2839
rect -2160 -2941 -2126 -2907
rect -2160 -3009 -2126 -2975
rect -2160 -3077 -2126 -3043
rect 2126 3043 2160 3077
rect 2126 2975 2160 3009
rect 2126 2907 2160 2941
rect 2126 2839 2160 2873
rect 2126 2771 2160 2805
rect 2126 2703 2160 2737
rect 2126 2635 2160 2669
rect 2126 2567 2160 2601
rect 2126 2499 2160 2533
rect 2126 2431 2160 2465
rect 2126 2363 2160 2397
rect 2126 2295 2160 2329
rect 2126 2227 2160 2261
rect 2126 2159 2160 2193
rect 2126 2091 2160 2125
rect 2126 2023 2160 2057
rect 2126 1955 2160 1989
rect 2126 1887 2160 1921
rect 2126 1819 2160 1853
rect 2126 1751 2160 1785
rect 2126 1683 2160 1717
rect 2126 1615 2160 1649
rect 2126 1547 2160 1581
rect 2126 1479 2160 1513
rect 2126 1411 2160 1445
rect 2126 1343 2160 1377
rect 2126 1275 2160 1309
rect 2126 1207 2160 1241
rect 2126 1139 2160 1173
rect 2126 1071 2160 1105
rect 2126 1003 2160 1037
rect 2126 935 2160 969
rect 2126 867 2160 901
rect 2126 799 2160 833
rect 2126 731 2160 765
rect 2126 663 2160 697
rect 2126 595 2160 629
rect 2126 527 2160 561
rect 2126 459 2160 493
rect 2126 391 2160 425
rect 2126 323 2160 357
rect 2126 255 2160 289
rect 2126 187 2160 221
rect 2126 119 2160 153
rect 2126 51 2160 85
rect 2126 -17 2160 17
rect 2126 -85 2160 -51
rect 2126 -153 2160 -119
rect 2126 -221 2160 -187
rect 2126 -289 2160 -255
rect 2126 -357 2160 -323
rect 2126 -425 2160 -391
rect 2126 -493 2160 -459
rect 2126 -561 2160 -527
rect 2126 -629 2160 -595
rect 2126 -697 2160 -663
rect 2126 -765 2160 -731
rect 2126 -833 2160 -799
rect 2126 -901 2160 -867
rect 2126 -969 2160 -935
rect 2126 -1037 2160 -1003
rect 2126 -1105 2160 -1071
rect 2126 -1173 2160 -1139
rect 2126 -1241 2160 -1207
rect 2126 -1309 2160 -1275
rect 2126 -1377 2160 -1343
rect 2126 -1445 2160 -1411
rect 2126 -1513 2160 -1479
rect 2126 -1581 2160 -1547
rect 2126 -1649 2160 -1615
rect 2126 -1717 2160 -1683
rect 2126 -1785 2160 -1751
rect 2126 -1853 2160 -1819
rect 2126 -1921 2160 -1887
rect 2126 -1989 2160 -1955
rect 2126 -2057 2160 -2023
rect 2126 -2125 2160 -2091
rect 2126 -2193 2160 -2159
rect 2126 -2261 2160 -2227
rect 2126 -2329 2160 -2295
rect 2126 -2397 2160 -2363
rect 2126 -2465 2160 -2431
rect 2126 -2533 2160 -2499
rect 2126 -2601 2160 -2567
rect 2126 -2669 2160 -2635
rect 2126 -2737 2160 -2703
rect 2126 -2805 2160 -2771
rect 2126 -2873 2160 -2839
rect 2126 -2941 2160 -2907
rect 2126 -3009 2160 -2975
rect -2160 -3145 -2126 -3111
rect 2126 -3077 2160 -3043
rect 2126 -3145 2160 -3111
rect -2160 -3213 -2126 -3179
rect 2126 -3213 2160 -3179
rect -2057 -3368 -2023 -3334
rect -1989 -3368 -1955 -3334
rect -1921 -3368 -1887 -3334
rect -1853 -3368 -1819 -3334
rect -1785 -3368 -1751 -3334
rect -1717 -3368 -1683 -3334
rect -1649 -3368 -1615 -3334
rect -1581 -3368 -1547 -3334
rect -1513 -3368 -1479 -3334
rect -1445 -3368 -1411 -3334
rect -1377 -3368 -1343 -3334
rect -1309 -3368 -1275 -3334
rect -1241 -3368 -1207 -3334
rect -1173 -3368 -1139 -3334
rect -1105 -3368 -1071 -3334
rect -1037 -3368 -1003 -3334
rect -969 -3368 -935 -3334
rect -901 -3368 -867 -3334
rect -833 -3368 -799 -3334
rect -765 -3368 -731 -3334
rect -697 -3368 -663 -3334
rect -629 -3368 -595 -3334
rect -561 -3368 -527 -3334
rect -493 -3368 -459 -3334
rect -425 -3368 -391 -3334
rect -357 -3368 -323 -3334
rect -289 -3368 -255 -3334
rect -221 -3368 -187 -3334
rect -153 -3368 -119 -3334
rect -85 -3368 -51 -3334
rect -17 -3368 17 -3334
rect 51 -3368 85 -3334
rect 119 -3368 153 -3334
rect 187 -3368 221 -3334
rect 255 -3368 289 -3334
rect 323 -3368 357 -3334
rect 391 -3368 425 -3334
rect 459 -3368 493 -3334
rect 527 -3368 561 -3334
rect 595 -3368 629 -3334
rect 663 -3368 697 -3334
rect 731 -3368 765 -3334
rect 799 -3368 833 -3334
rect 867 -3368 901 -3334
rect 935 -3368 969 -3334
rect 1003 -3368 1037 -3334
rect 1071 -3368 1105 -3334
rect 1139 -3368 1173 -3334
rect 1207 -3368 1241 -3334
rect 1275 -3368 1309 -3334
rect 1343 -3368 1377 -3334
rect 1411 -3368 1445 -3334
rect 1479 -3368 1513 -3334
rect 1547 -3368 1581 -3334
rect 1615 -3368 1649 -3334
rect 1683 -3368 1717 -3334
rect 1751 -3368 1785 -3334
rect 1819 -3368 1853 -3334
rect 1887 -3368 1921 -3334
rect 1955 -3368 1989 -3334
rect 2023 -3368 2057 -3334
<< locali >>
rect -2160 3334 -2057 3368
rect -2023 3334 -1989 3368
rect -1955 3334 -1921 3368
rect -1887 3334 -1853 3368
rect -1819 3334 -1785 3368
rect -1751 3334 -1717 3368
rect -1683 3334 -1649 3368
rect -1615 3334 -1581 3368
rect -1547 3334 -1513 3368
rect -1479 3334 -1445 3368
rect -1411 3334 -1377 3368
rect -1343 3334 -1309 3368
rect -1275 3334 -1241 3368
rect -1207 3334 -1173 3368
rect -1139 3334 -1105 3368
rect -1071 3334 -1037 3368
rect -1003 3334 -969 3368
rect -935 3334 -901 3368
rect -867 3334 -833 3368
rect -799 3334 -765 3368
rect -731 3334 -697 3368
rect -663 3334 -629 3368
rect -595 3334 -561 3368
rect -527 3334 -493 3368
rect -459 3334 -425 3368
rect -391 3334 -357 3368
rect -323 3334 -289 3368
rect -255 3334 -221 3368
rect -187 3334 -153 3368
rect -119 3334 -85 3368
rect -51 3334 -17 3368
rect 17 3334 51 3368
rect 85 3334 119 3368
rect 153 3334 187 3368
rect 221 3334 255 3368
rect 289 3334 323 3368
rect 357 3334 391 3368
rect 425 3334 459 3368
rect 493 3334 527 3368
rect 561 3334 595 3368
rect 629 3334 663 3368
rect 697 3334 731 3368
rect 765 3334 799 3368
rect 833 3334 867 3368
rect 901 3334 935 3368
rect 969 3334 1003 3368
rect 1037 3334 1071 3368
rect 1105 3334 1139 3368
rect 1173 3334 1207 3368
rect 1241 3334 1275 3368
rect 1309 3334 1343 3368
rect 1377 3334 1411 3368
rect 1445 3334 1479 3368
rect 1513 3334 1547 3368
rect 1581 3334 1615 3368
rect 1649 3334 1683 3368
rect 1717 3334 1751 3368
rect 1785 3334 1819 3368
rect 1853 3334 1887 3368
rect 1921 3334 1955 3368
rect 1989 3334 2023 3368
rect 2057 3334 2160 3368
rect -2160 3213 -2126 3334
rect -2160 3145 -2126 3179
rect 2126 3213 2160 3334
rect -2160 3077 -2126 3111
rect -1952 3154 1952 3156
rect -1952 3110 -1921 3154
rect 1921 3110 1952 3154
rect -1952 3076 -1925 3110
rect 1925 3076 1952 3110
rect -1952 3052 -1921 3076
rect 1921 3052 1952 3076
rect -1952 3050 1952 3052
rect 2126 3145 2160 3179
rect 2126 3077 2160 3111
rect -2160 3009 -2126 3043
rect -2160 2941 -2126 2975
rect -2160 2873 -2126 2907
rect -2160 2805 -2126 2839
rect -2160 2737 -2126 2771
rect -2160 2669 -2126 2703
rect -2160 2601 -2126 2635
rect -2160 2533 -2126 2567
rect -2160 2465 -2126 2499
rect -2160 2397 -2126 2431
rect -2160 2329 -2126 2363
rect -2160 2261 -2126 2295
rect -2160 2193 -2126 2227
rect -2160 2125 -2126 2159
rect -2160 2057 -2126 2091
rect -2160 1989 -2126 2023
rect -2160 1921 -2126 1955
rect -2160 1853 -2126 1887
rect -2160 1785 -2126 1819
rect -2160 1717 -2126 1751
rect -2160 1649 -2126 1683
rect -2160 1581 -2126 1615
rect -2160 1513 -2126 1547
rect -2160 1445 -2126 1479
rect -2160 1377 -2126 1411
rect -2160 1309 -2126 1343
rect -2160 1241 -2126 1275
rect -2160 1173 -2126 1207
rect -2160 1105 -2126 1139
rect -2160 1037 -2126 1071
rect -2160 969 -2126 1003
rect -2160 901 -2126 935
rect -2160 833 -2126 867
rect -2160 765 -2126 799
rect -2160 697 -2126 731
rect -2160 629 -2126 663
rect -2160 561 -2126 595
rect -2160 493 -2126 527
rect -2160 425 -2126 459
rect -2160 357 -2126 391
rect -2160 289 -2126 323
rect -2160 221 -2126 255
rect -2160 153 -2126 187
rect -2160 85 -2126 119
rect -2160 17 -2126 51
rect -2160 -51 -2126 -17
rect -2160 -119 -2126 -85
rect -2160 -187 -2126 -153
rect -2160 -255 -2126 -221
rect -2160 -323 -2126 -289
rect -2160 -391 -2126 -357
rect -2160 -459 -2126 -425
rect -2160 -527 -2126 -493
rect -2160 -595 -2126 -561
rect -2160 -663 -2126 -629
rect -2160 -731 -2126 -697
rect -2160 -799 -2126 -765
rect -2160 -867 -2126 -833
rect -2160 -935 -2126 -901
rect -2160 -1003 -2126 -969
rect -2160 -1071 -2126 -1037
rect -2160 -1139 -2126 -1105
rect -2160 -1207 -2126 -1173
rect -2160 -1275 -2126 -1241
rect -2160 -1343 -2126 -1309
rect -2160 -1411 -2126 -1377
rect -2160 -1479 -2126 -1445
rect -2160 -1547 -2126 -1513
rect -2160 -1615 -2126 -1581
rect -2160 -1683 -2126 -1649
rect -2160 -1751 -2126 -1717
rect -2160 -1819 -2126 -1785
rect -2160 -1887 -2126 -1853
rect -2160 -1955 -2126 -1921
rect -2160 -2023 -2126 -1989
rect -2160 -2091 -2126 -2057
rect -2160 -2159 -2126 -2125
rect -2160 -2227 -2126 -2193
rect -2160 -2295 -2126 -2261
rect -2160 -2363 -2126 -2329
rect -2160 -2431 -2126 -2397
rect -2160 -2499 -2126 -2465
rect -2160 -2567 -2126 -2533
rect -2160 -2635 -2126 -2601
rect -2160 -2703 -2126 -2669
rect -2160 -2771 -2126 -2737
rect -2160 -2839 -2126 -2805
rect -2160 -2907 -2126 -2873
rect -2160 -2975 -2126 -2941
rect -2160 -3043 -2126 -3009
rect 2126 3009 2160 3043
rect 2126 2941 2160 2975
rect 2126 2873 2160 2907
rect 2126 2805 2160 2839
rect 2126 2737 2160 2771
rect 2126 2669 2160 2703
rect 2126 2601 2160 2635
rect 2126 2533 2160 2567
rect 2126 2465 2160 2499
rect 2126 2397 2160 2431
rect 2126 2329 2160 2363
rect 2126 2261 2160 2295
rect 2126 2193 2160 2227
rect 2126 2125 2160 2159
rect 2126 2057 2160 2091
rect 2126 1989 2160 2023
rect 2126 1921 2160 1955
rect 2126 1853 2160 1887
rect 2126 1785 2160 1819
rect 2126 1717 2160 1751
rect 2126 1649 2160 1683
rect 2126 1581 2160 1615
rect 2126 1513 2160 1547
rect 2126 1445 2160 1479
rect 2126 1377 2160 1411
rect 2126 1309 2160 1343
rect 2126 1241 2160 1275
rect 2126 1173 2160 1207
rect 2126 1105 2160 1139
rect 2126 1037 2160 1071
rect 2126 969 2160 1003
rect 2126 901 2160 935
rect 2126 833 2160 867
rect 2126 765 2160 799
rect 2126 697 2160 731
rect 2126 629 2160 663
rect 2126 561 2160 595
rect 2126 493 2160 527
rect 2126 425 2160 459
rect 2126 357 2160 391
rect 2126 289 2160 323
rect 2126 221 2160 255
rect 2126 153 2160 187
rect 2126 85 2160 119
rect 2126 17 2160 51
rect 2126 -51 2160 -17
rect 2126 -119 2160 -85
rect 2126 -187 2160 -153
rect 2126 -255 2160 -221
rect 2126 -323 2160 -289
rect 2126 -391 2160 -357
rect 2126 -459 2160 -425
rect 2126 -527 2160 -493
rect 2126 -595 2160 -561
rect 2126 -663 2160 -629
rect 2126 -731 2160 -697
rect 2126 -799 2160 -765
rect 2126 -867 2160 -833
rect 2126 -935 2160 -901
rect 2126 -1003 2160 -969
rect 2126 -1071 2160 -1037
rect 2126 -1139 2160 -1105
rect 2126 -1207 2160 -1173
rect 2126 -1275 2160 -1241
rect 2126 -1343 2160 -1309
rect 2126 -1411 2160 -1377
rect 2126 -1479 2160 -1445
rect 2126 -1547 2160 -1513
rect 2126 -1615 2160 -1581
rect 2126 -1683 2160 -1649
rect 2126 -1751 2160 -1717
rect 2126 -1819 2160 -1785
rect 2126 -1887 2160 -1853
rect 2126 -1955 2160 -1921
rect 2126 -2023 2160 -1989
rect 2126 -2091 2160 -2057
rect 2126 -2159 2160 -2125
rect 2126 -2227 2160 -2193
rect 2126 -2295 2160 -2261
rect 2126 -2363 2160 -2329
rect 2126 -2431 2160 -2397
rect 2126 -2499 2160 -2465
rect 2126 -2567 2160 -2533
rect 2126 -2635 2160 -2601
rect 2126 -2703 2160 -2669
rect 2126 -2771 2160 -2737
rect 2126 -2839 2160 -2805
rect 2126 -2907 2160 -2873
rect 2126 -2975 2160 -2941
rect 2126 -3043 2160 -3009
rect -2160 -3111 -2126 -3077
rect -2160 -3179 -2126 -3145
rect -1952 -3052 1952 -3050
rect -1952 -3076 -1921 -3052
rect 1921 -3076 1952 -3052
rect -1952 -3110 -1925 -3076
rect 1925 -3110 1952 -3076
rect -1952 -3154 -1921 -3110
rect 1921 -3154 1952 -3110
rect -1952 -3156 1952 -3154
rect 2126 -3111 2160 -3077
rect -2160 -3334 -2126 -3213
rect 2126 -3179 2160 -3145
rect 2126 -3334 2160 -3213
rect -2160 -3368 -2057 -3334
rect -2023 -3368 -1989 -3334
rect -1955 -3368 -1921 -3334
rect -1887 -3368 -1853 -3334
rect -1819 -3368 -1785 -3334
rect -1751 -3368 -1717 -3334
rect -1683 -3368 -1649 -3334
rect -1615 -3368 -1581 -3334
rect -1547 -3368 -1513 -3334
rect -1479 -3368 -1445 -3334
rect -1411 -3368 -1377 -3334
rect -1343 -3368 -1309 -3334
rect -1275 -3368 -1241 -3334
rect -1207 -3368 -1173 -3334
rect -1139 -3368 -1105 -3334
rect -1071 -3368 -1037 -3334
rect -1003 -3368 -969 -3334
rect -935 -3368 -901 -3334
rect -867 -3368 -833 -3334
rect -799 -3368 -765 -3334
rect -731 -3368 -697 -3334
rect -663 -3368 -629 -3334
rect -595 -3368 -561 -3334
rect -527 -3368 -493 -3334
rect -459 -3368 -425 -3334
rect -391 -3368 -357 -3334
rect -323 -3368 -289 -3334
rect -255 -3368 -221 -3334
rect -187 -3368 -153 -3334
rect -119 -3368 -85 -3334
rect -51 -3368 -17 -3334
rect 17 -3368 51 -3334
rect 85 -3368 119 -3334
rect 153 -3368 187 -3334
rect 221 -3368 255 -3334
rect 289 -3368 323 -3334
rect 357 -3368 391 -3334
rect 425 -3368 459 -3334
rect 493 -3368 527 -3334
rect 561 -3368 595 -3334
rect 629 -3368 663 -3334
rect 697 -3368 731 -3334
rect 765 -3368 799 -3334
rect 833 -3368 867 -3334
rect 901 -3368 935 -3334
rect 969 -3368 1003 -3334
rect 1037 -3368 1071 -3334
rect 1105 -3368 1139 -3334
rect 1173 -3368 1207 -3334
rect 1241 -3368 1275 -3334
rect 1309 -3368 1343 -3334
rect 1377 -3368 1411 -3334
rect 1445 -3368 1479 -3334
rect 1513 -3368 1547 -3334
rect 1581 -3368 1615 -3334
rect 1649 -3368 1683 -3334
rect 1717 -3368 1751 -3334
rect 1785 -3368 1819 -3334
rect 1853 -3368 1887 -3334
rect 1921 -3368 1955 -3334
rect 1989 -3368 2023 -3334
rect 2057 -3368 2160 -3334
<< viali >>
rect -1925 3076 -1921 3110
rect -1921 3076 -1891 3110
rect -1853 3076 -1819 3110
rect -1781 3076 -1747 3110
rect -1709 3076 -1675 3110
rect -1637 3076 -1603 3110
rect -1565 3076 -1531 3110
rect -1493 3076 -1459 3110
rect -1421 3076 -1387 3110
rect -1349 3076 -1315 3110
rect -1277 3076 -1243 3110
rect -1205 3076 -1171 3110
rect -1133 3076 -1099 3110
rect -1061 3076 -1027 3110
rect -989 3076 -955 3110
rect -917 3076 -883 3110
rect -845 3076 -811 3110
rect -773 3076 -739 3110
rect -701 3076 -667 3110
rect -629 3076 -595 3110
rect -557 3076 -523 3110
rect -485 3076 -451 3110
rect -413 3076 -379 3110
rect -341 3076 -307 3110
rect -269 3076 -235 3110
rect -197 3076 -163 3110
rect -125 3076 -91 3110
rect -53 3076 -19 3110
rect 19 3076 53 3110
rect 91 3076 125 3110
rect 163 3076 197 3110
rect 235 3076 269 3110
rect 307 3076 341 3110
rect 379 3076 413 3110
rect 451 3076 485 3110
rect 523 3076 557 3110
rect 595 3076 629 3110
rect 667 3076 701 3110
rect 739 3076 773 3110
rect 811 3076 845 3110
rect 883 3076 917 3110
rect 955 3076 989 3110
rect 1027 3076 1061 3110
rect 1099 3076 1133 3110
rect 1171 3076 1205 3110
rect 1243 3076 1277 3110
rect 1315 3076 1349 3110
rect 1387 3076 1421 3110
rect 1459 3076 1493 3110
rect 1531 3076 1565 3110
rect 1603 3076 1637 3110
rect 1675 3076 1709 3110
rect 1747 3076 1781 3110
rect 1819 3076 1853 3110
rect 1891 3076 1921 3110
rect 1921 3076 1925 3110
rect -1925 -3110 -1921 -3076
rect -1921 -3110 -1891 -3076
rect -1853 -3110 -1819 -3076
rect -1781 -3110 -1747 -3076
rect -1709 -3110 -1675 -3076
rect -1637 -3110 -1603 -3076
rect -1565 -3110 -1531 -3076
rect -1493 -3110 -1459 -3076
rect -1421 -3110 -1387 -3076
rect -1349 -3110 -1315 -3076
rect -1277 -3110 -1243 -3076
rect -1205 -3110 -1171 -3076
rect -1133 -3110 -1099 -3076
rect -1061 -3110 -1027 -3076
rect -989 -3110 -955 -3076
rect -917 -3110 -883 -3076
rect -845 -3110 -811 -3076
rect -773 -3110 -739 -3076
rect -701 -3110 -667 -3076
rect -629 -3110 -595 -3076
rect -557 -3110 -523 -3076
rect -485 -3110 -451 -3076
rect -413 -3110 -379 -3076
rect -341 -3110 -307 -3076
rect -269 -3110 -235 -3076
rect -197 -3110 -163 -3076
rect -125 -3110 -91 -3076
rect -53 -3110 -19 -3076
rect 19 -3110 53 -3076
rect 91 -3110 125 -3076
rect 163 -3110 197 -3076
rect 235 -3110 269 -3076
rect 307 -3110 341 -3076
rect 379 -3110 413 -3076
rect 451 -3110 485 -3076
rect 523 -3110 557 -3076
rect 595 -3110 629 -3076
rect 667 -3110 701 -3076
rect 739 -3110 773 -3076
rect 811 -3110 845 -3076
rect 883 -3110 917 -3076
rect 955 -3110 989 -3076
rect 1027 -3110 1061 -3076
rect 1099 -3110 1133 -3076
rect 1171 -3110 1205 -3076
rect 1243 -3110 1277 -3076
rect 1315 -3110 1349 -3076
rect 1387 -3110 1421 -3076
rect 1459 -3110 1493 -3076
rect 1531 -3110 1565 -3076
rect 1603 -3110 1637 -3076
rect 1675 -3110 1709 -3076
rect 1747 -3110 1781 -3076
rect 1819 -3110 1853 -3076
rect 1891 -3110 1921 -3076
rect 1921 -3110 1925 -3076
<< metal1 >>
rect -1960 3110 1960 3126
rect -1960 3076 -1925 3110
rect -1891 3076 -1853 3110
rect -1819 3076 -1781 3110
rect -1747 3076 -1709 3110
rect -1675 3076 -1637 3110
rect -1603 3076 -1565 3110
rect -1531 3076 -1493 3110
rect -1459 3076 -1421 3110
rect -1387 3076 -1349 3110
rect -1315 3076 -1277 3110
rect -1243 3076 -1205 3110
rect -1171 3076 -1133 3110
rect -1099 3076 -1061 3110
rect -1027 3076 -989 3110
rect -955 3076 -917 3110
rect -883 3076 -845 3110
rect -811 3076 -773 3110
rect -739 3076 -701 3110
rect -667 3076 -629 3110
rect -595 3076 -557 3110
rect -523 3076 -485 3110
rect -451 3076 -413 3110
rect -379 3076 -341 3110
rect -307 3076 -269 3110
rect -235 3076 -197 3110
rect -163 3076 -125 3110
rect -91 3076 -53 3110
rect -19 3076 19 3110
rect 53 3076 91 3110
rect 125 3076 163 3110
rect 197 3076 235 3110
rect 269 3076 307 3110
rect 341 3076 379 3110
rect 413 3076 451 3110
rect 485 3076 523 3110
rect 557 3076 595 3110
rect 629 3076 667 3110
rect 701 3076 739 3110
rect 773 3076 811 3110
rect 845 3076 883 3110
rect 917 3076 955 3110
rect 989 3076 1027 3110
rect 1061 3076 1099 3110
rect 1133 3076 1171 3110
rect 1205 3076 1243 3110
rect 1277 3076 1315 3110
rect 1349 3076 1387 3110
rect 1421 3076 1459 3110
rect 1493 3076 1531 3110
rect 1565 3076 1603 3110
rect 1637 3076 1675 3110
rect 1709 3076 1747 3110
rect 1781 3076 1819 3110
rect 1853 3076 1891 3110
rect 1925 3076 1960 3110
rect -1960 3061 1960 3076
rect -1960 -3076 1960 -3061
rect -1960 -3110 -1925 -3076
rect -1891 -3110 -1853 -3076
rect -1819 -3110 -1781 -3076
rect -1747 -3110 -1709 -3076
rect -1675 -3110 -1637 -3076
rect -1603 -3110 -1565 -3076
rect -1531 -3110 -1493 -3076
rect -1459 -3110 -1421 -3076
rect -1387 -3110 -1349 -3076
rect -1315 -3110 -1277 -3076
rect -1243 -3110 -1205 -3076
rect -1171 -3110 -1133 -3076
rect -1099 -3110 -1061 -3076
rect -1027 -3110 -989 -3076
rect -955 -3110 -917 -3076
rect -883 -3110 -845 -3076
rect -811 -3110 -773 -3076
rect -739 -3110 -701 -3076
rect -667 -3110 -629 -3076
rect -595 -3110 -557 -3076
rect -523 -3110 -485 -3076
rect -451 -3110 -413 -3076
rect -379 -3110 -341 -3076
rect -307 -3110 -269 -3076
rect -235 -3110 -197 -3076
rect -163 -3110 -125 -3076
rect -91 -3110 -53 -3076
rect -19 -3110 19 -3076
rect 53 -3110 91 -3076
rect 125 -3110 163 -3076
rect 197 -3110 235 -3076
rect 269 -3110 307 -3076
rect 341 -3110 379 -3076
rect 413 -3110 451 -3076
rect 485 -3110 523 -3076
rect 557 -3110 595 -3076
rect 629 -3110 667 -3076
rect 701 -3110 739 -3076
rect 773 -3110 811 -3076
rect 845 -3110 883 -3076
rect 917 -3110 955 -3076
rect 989 -3110 1027 -3076
rect 1061 -3110 1099 -3076
rect 1133 -3110 1171 -3076
rect 1205 -3110 1243 -3076
rect 1277 -3110 1315 -3076
rect 1349 -3110 1387 -3076
rect 1421 -3110 1459 -3076
rect 1493 -3110 1531 -3076
rect 1565 -3110 1603 -3076
rect 1637 -3110 1675 -3076
rect 1709 -3110 1747 -3076
rect 1781 -3110 1819 -3076
rect 1853 -3110 1891 -3076
rect 1925 -3110 1960 -3076
rect -1960 -3126 1960 -3110
<< end >>
