magic
tech sky130A
magscale 1 2
timestamp 1713591521
<< error_p >>
rect 0 284 1922 320
<< metal4 >>
rect 0 260 1922 284
rect 0 24 43 260
rect 279 24 363 260
rect 599 24 683 260
rect 919 24 1003 260
rect 1239 24 1323 260
rect 1559 24 1643 260
rect 1879 24 1922 260
rect 0 0 1922 24
<< via4 >>
rect 43 24 279 260
rect 363 24 599 260
rect 683 24 919 260
rect 1003 24 1239 260
rect 1323 24 1559 260
rect 1643 24 1879 260
<< metal5 >>
rect 0 260 1922 284
rect 0 24 43 260
rect 279 24 363 260
rect 599 24 683 260
rect 919 24 1003 260
rect 1239 24 1323 260
rect 1559 24 1643 260
rect 1879 24 1922 260
rect 0 0 1922 24
<< end >>
