* NGSPICE file created from ONES_COUNTER_pex.ext - technology: sky130A

.subckt ONES_COUNTER_pex VGND VPWR clk rst pulse ready ones[0] ones[1] ones[2] ones[3] ones[4] ones[5]
+ ones[6] ones[7] ones[8] ones[9] ones[10]
X0 a_4414_4399# counter\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.17515 ps=1.265 w=0.42 l=0.15
X1 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=142.45384 ps=1.33502k w=0.87 l=1.97
X2 a_8268_2741# net6 a_8397_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3 _081_ net3 a_5446_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
X4 a_1932_10933# _023_ a_1860_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X5 a_2419_2767# _045_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.15 ps=1.3 w=1 l=0.15
X6 VPWR counter\[4\] a_3847_6727# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X7 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X8 a_4135_4373# counter\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_4616_4399# counter\[1\] a_4510_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0798 ps=0.8 w=0.42 l=0.15
X10 VGND net10 a_9043_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X11 VGND a_3099_9117# a_3267_9019# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X12 a_9079_6031# a_8381_6037# a_8822_6005# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X13 VGND _069_ _006_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND a_7102_6575# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X15 VGND a_5433_7637# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X16 VPWR _075_ a_10103_9991# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X17 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=90.401054 ps=954.98 w=0.55 l=2.89
X18 a_3965_8751# a_3799_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_8017_4943# _002_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X20 _072_ a_10134_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X21 a_7996_9001# counter\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X22 a_6541_8213# a_6375_8213# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 VPWR a_10103_9514# _013_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X24 a_10337_9839# _075_ a_10265_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X25 a_7263_7637# net6 a_7744_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X26 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X27 VGND net1 a_9926_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X28 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X29 VPWR clknet_1_1__leaf_clk a_6743_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X30 a_1915_5639# a_2011_5461# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X31 a_5437_4399# a_5271_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X32 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X33 VPWR _043_ a_2790_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.18 ps=1.36 w=1 l=0.15
X34 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X35 a_8293_5487# net6 a_8205_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X36 VGND net3 a_8399_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X37 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X38 a_2668_4405# _024_ a_2596_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X39 a_7843_5737# _061_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X40 a_9411_7119# net2 _052_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.175 ps=1.35 w=1 l=0.15
X41 ones[0] a_9779_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X42 a_9117_7663# a_8951_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X43 a_9735_5639# net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.134875 ps=1.065 w=0.65 l=0.15
X44 VPWR _024_ a_2787_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X45 clknet_0_clk a_5433_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X46 VPWR a_3847_3463# _033_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X47 a_10199_3285# pulse VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X48 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X49 a_2325_5263# counter\[9\] a_2229_5263# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X50 a_2941_6351# _047_ a_2869_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.06825 ps=0.86 w=0.65 l=0.15
X51 VPWR counter\[7\] _076_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X52 counter\[8\] a_7407_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X53 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X54 VGND counter\[0\] a_5018_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X55 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X56 VPWR a_9815_8029# a_9983_7931# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X57 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X58 a_10199_2197# rst VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X59 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X60 VPWR a_4227_9513# a_4234_9417# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X61 a_9079_6031# a_8215_6037# a_8822_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X62 VGND a_8367_7337# a_8374_7241# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X63 a_6324_10029# _064_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X64 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X65 VPWR a_3099_9117# a_3267_9019# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X66 a_8767_10749# counter\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X67 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X68 clknet_1_0__leaf_clk a_3593_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X69 a_3965_7125# a_3799_7125# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X70 VPWR net9 a_9739_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X71 a_7323_8207# a_6541_8213# a_7239_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X72 a_9117_6575# a_8951_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X73 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X74 _068_ a_8767_10749# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X75 VPWR a_7102_6575# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X76 a_2593_2223# _053_ a_2511_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X77 VPWR a_3593_8181# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X78 VGND a_4406_7093# a_4364_7497# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X79 VPWR a_4491_6263# _057_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X80 VPWR counter\[8\] a_3476_7351# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1087 ps=1.36 w=0.42 l=0.15
X81 _012_ _085_ a_1505_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X82 VGND a_8268_2741# _023_ VGND sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X83 a_9558_6687# a_9390_6941# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X84 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X85 a_8355_4074# _048_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X86 a_7987_7351# a_8083_7351# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X87 VGND a_9815_8029# a_9983_7931# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X88 VGND net12 _044_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X89 VPWR a_8075_3285# a_7711_3463# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X90 VPWR clknet_1_1__leaf_clk a_6375_8213# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X91 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X92 VPWR net14 _080_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X93 VPWR net14 a_9963_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X94 a_5496_9269# _024_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.101875 ps=0.99 w=0.42 l=0.15
X95 VPWR _053_ a_6835_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X96 VGND counter\[2\] a_9122_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X97 VGND a_4894_6549# a_4823_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X98 a_4798_5737# a_5018_5461# _050_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X99 a_6612_3829# _068_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X100 a_7343_7351# a_7616_7351# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1085 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X101 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X102 a_8397_3087# _083_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X103 a_1915_5639# a_2011_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X104 a_5625_4399# _016_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X105 a_4406_8863# a_4238_9117# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X106 _024_ net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X107 VPWR a_9247_6005# a_9163_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X108 VPWR clknet_1_0__leaf_clk a_3799_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X109 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X110 VPWR net2 a_2971_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X111 _014_ a_2776_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X112 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X113 a_9815_6941# a_9117_6575# a_9558_6687# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X114 VGND a_3819_4917# net3 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X115 _058_ counter\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X116 a_1559_2473# counter\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X117 a_9739_6005# _028_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.31245 ps=1.68 w=0.42 l=0.15
X118 _000_ a_2879_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X119 VPWR a_5050_4917# a_4977_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X120 VPWR _033_ a_5271_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X121 VGND a_5043_4564# _015_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X122 a_7515_6031# a_6651_6037# a_7258_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X123 a_2409_4445# _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X124 VGND a_5475_4917# a_5433_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X125 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X126 a_4153_7119# _015_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X128 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X129 VPWR a_6979_10901# _007_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X131 VGND a_9735_5639# _085_ VGND sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
X132 a_9117_6575# a_8951_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X133 a_9815_6941# a_8951_6575# a_9558_6687# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X134 VGND clknet_1_0__leaf_clk a_3799_7125# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X135 a_5513_10089# counter\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X136 a_8921_7497# a_8374_7241# a_8574_7396# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X137 net11 a_9983_6843# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X138 VPWR a_7711_3463# _051_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X139 a_2676_2767# _039_ a_2419_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.1375 ps=1.275 w=1 l=0.15
X140 a_4609_4949# a_4443_4949# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X141 a_3847_9527# a_3943_9527# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X142 _083_ a_9926_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X143 a_2787_6031# _047_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.15 ps=1.3 w=1 l=0.15
X144 a_6324_10029# _064_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.101875 ps=0.99 w=0.42 l=0.15
X145 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X146 VPWR net9 a_10239_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X147 VGND net12 a_6060_6549# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X148 clknet_1_0__leaf_clk a_3593_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X149 VGND a_3300_9269# _053_ VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X150 VPWR a_1915_5639# counter\[10\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X151 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X152 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X153 VGND _057_ a_1775_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X154 a_3521_3971# _053_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X155 a_4143_6397# _086_ a_4047_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X156 _020_ a_2419_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3125 ps=1.625 w=1 l=0.15
X157 a_9868_5487# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.112125 ps=0.995 w=0.65 l=0.15
X158 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X159 _059_ a_9122_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X160 VPWR net12 _040_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X161 VGND a_5433_7637# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X162 VPWR _080_ a_5363_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.265 ps=2.53 w=1 l=0.15
X163 a_3867_9813# a_4035_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X164 a_10103_9991# _076_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X165 VGND a_10103_9514# _013_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X166 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X167 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X168 a_2849_5487# a_2295_5461# a_2502_5461# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X169 VGND a_7531_2741# _047_ VGND sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X170 VGND _033_ a_5271_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X171 VPWR a_7683_6005# a_7599_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X172 net11 a_9983_6843# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X173 VPWR _069_ a_1559_2473# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X174 VPWR a_3593_8181# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X175 a_9201_4399# net11 a_9117_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X176 VPWR _054_ a_2879_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X177 a_7090_6031# a_6651_6037# a_7005_6031# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X178 a_4403_6549# a_4687_6549# a_4622_6575# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X179 a_4663_9117# a_3799_8751# a_4406_8863# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X180 a_2401_8751# a_2235_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X181 a_8265_10721# net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X182 a_2678_5853# a_2431_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X183 VPWR a_9983_6843# a_9899_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X184 a_2401_7663# a_2235_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X186 a_2511_2223# _058_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X187 a_8863_8527# _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.105625 ps=0.975 w=0.65 l=0.15
X188 VGND a_6303_4667# a_6261_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X189 VPWR net13 a_7749_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X190 a_4491_6263# _053_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X191 clknet_1_1__leaf_clk a_7102_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X192 a_3847_6727# counter\[5\] a_4081_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X193 VGND a_5433_7637# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X194 a_5613_7439# counter\[9\] a_5529_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X195 a_2007_7828# _042_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X196 a_4406_8863# a_4238_9117# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X197 a_2589_7663# _004_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X198 VGND a_4589_3829# _029_ VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X199 VPWR a_5433_7637# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X200 a_4491_6263# _053_ a_4725_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X201 VGND a_3847_6727# _065_ VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X203 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X204 VPWR _053_ a_10136_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.195 ps=1.39 w=1 l=0.15
X205 _075_ a_1465_2473# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X207 a_9815_8029# a_8951_7663# a_9558_7775# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X208 a_10134_10927# counter\[8\] a_9965_11177# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X209 _002_ a_6375_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X210 a_3203_7351# a_3476_7351# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1085 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X211 a_6093_8527# counter\[8\] a_5997_8527# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X212 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X213 a_7216_6409# a_6817_6037# a_7090_6031# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X214 VGND net9 a_10239_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X215 VGND a_6579_9019# counter\[1\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X216 a_4511_3087# _080_ a_4415_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X217 a_8013_3087# net11 a_7917_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X218 counter\[8\] a_7407_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X219 VGND a_3593_8181# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X221 a_3847_3463# a_4120_3291# a_4078_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.107825 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X222 VGND a_7987_7351# net6 VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X223 _080_ net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X225 a_1489_4649# counter\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X226 VPWR _083_ a_4807_3855# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X227 VGND _037_ a_2668_4405# VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X228 a_6537_8751# a_5547_8751# a_6411_9117# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X229 a_8803_9295# a_8105_9301# a_8546_9269# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X230 VGND net4 _046_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X231 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X232 a_7845_3311# counter\[4\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X233 VPWR clknet_0_clk a_7102_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X234 clknet_0_clk a_5433_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X235 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X236 VPWR a_4831_9019# a_4747_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X237 a_2849_5487# a_2302_5761# a_2502_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X238 a_2230_5487# a_1915_5639# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X239 VGND a_1915_5639# counter\[10\] VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X240 a_8945_8207# _078_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X241 a_4702_10205# a_4455_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X242 VGND a_8091_10615# _034_ VGND sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X243 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X244 a_9011_3285# net8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.0777 ps=0.79 w=0.42 l=0.15
X245 VGND a_6579_9019# a_6537_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X246 a_8123_5487# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X247 a_7729_10927# _031_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X248 VGND net5 a_9503_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X249 _005_ a_5823_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X250 VPWR counter\[10\] _078_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X251 VPWR net3 a_9779_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X252 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X253 _024_ net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X254 VPWR a_9983_7931# a_9899_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X255 ones[0] a_9779_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X256 VPWR net7 a_9011_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X257 VGND a_3394_4917# a_3352_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X258 VGND a_2842_7775# a_2800_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X259 a_8105_9301# a_7939_9301# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X260 VPWR clknet_1_1__leaf_clk a_7663_4949# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X261 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X262 a_4526_9813# a_4319_9813# a_4702_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X263 a_10136_4943# _061_ a_10045_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1525 ps=1.305 w=1 l=0.15
X264 a_4455_9839# a_4319_9813# a_4035_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X265 VPWR a_9011_3285# _031_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.165 ps=1.33 w=1 l=0.15
X266 a_3513_6825# _070_ _006_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X267 _048_ a_3137_4765# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X268 _053_ a_3300_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X269 a_2842_8863# a_2674_9117# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X270 a_6099_10089# counter\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X271 VPWR a_6579_9019# counter\[1\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X272 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X273 _086_ a_7263_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X275 a_4981_6263# _036_ a_5144_6147# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X276 a_7625_5461# counter\[5\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X277 VGND net1 a_4511_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X278 a_4747_8029# a_3965_7663# a_4663_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X279 a_1673_10973# _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X280 VGND a_3651_4943# a_3819_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X282 VPWR _053_ _070_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X283 a_8325_7119# a_7987_7351# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X284 VGND a_6612_3829# _069_ VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X286 VPWR a_6135_4765# a_6303_4667# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X288 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X289 counter\[5\] a_7775_4667# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X290 VGND clk a_5433_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X291 a_9551_9527# net8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X293 a_6335_5461# _053_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X294 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X295 a_7987_7828# _077_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X296 a_4254_9839# a_3867_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X297 VPWR a_5878_4511# a_5805_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X298 _082_ a_4225_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X299 VGND counter\[10\] a_2409_5263# VGND sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.183625 ps=1.215 w=0.65 l=0.15
X300 counter\[6\] a_5475_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X301 VPWR counter\[1\] a_4351_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X302 a_4434_9572# a_4227_9513# a_4610_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X303 a_2397_9839# a_1407_9839# a_2271_10205# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X304 a_9661_7439# _049_ _052_ VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.169 ps=1.82 w=0.65 l=0.15
X305 a_3141_4943# _011_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X307 a_2589_7663# _004_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X308 clknet_0_clk a_5433_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X309 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X310 VGND a_2439_10107# a_2397_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X311 a_5805_4765# a_5271_4399# a_5710_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X312 VGND a_6135_4765# a_6303_4667# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X313 a_4610_9295# a_4363_9673# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X314 a_9713_9661# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X315 VPWR a_1761_2999# _032_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X316 VPWR clknet_1_0__leaf_clk a_2235_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X317 VGND _081_ _011_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X318 a_8355_4074# _048_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X319 a_8503_7497# a_8367_7337# a_8083_7351# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X320 clknet_1_0__leaf_clk a_3593_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X321 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X322 _067_ a_3521_3971# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X323 clknet_1_0__leaf_clk a_3593_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X324 a_8381_6037# a_8215_6037# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X325 a_8378_9295# a_7939_9301# a_8293_9295# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X326 a_4434_9572# a_4234_9417# a_4583_9661# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X327 a_2011_5461# a_2295_5461# a_2230_5487# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X328 a_4747_7119# a_3965_7125# a_4663_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X329 _025_ a_1773_11191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X330 a_7711_3463# a_8075_3285# a_8033_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X331 a_2007_7828# _042_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X332 a_2665_2223# _058_ a_2593_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X333 VPWR a_7102_6575# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X334 a_9290_3311# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.17515 ps=1.265 w=0.42 l=0.15
X335 a_7365_8585# a_6375_8213# a_7239_8207# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X336 a_3225_8751# a_2235_8751# a_3099_9117# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X337 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X338 a_8887_9295# a_8105_9301# a_8803_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X339 a_5356_9615# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X340 a_9492_3311# net8 a_9386_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0798 ps=0.8 w=0.42 l=0.15
X341 VPWR net3 a_4621_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X342 a_4135_4373# counter\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.27995 ps=1.615 w=0.42 l=0.15
X343 a_3158_6031# _043_ a_3044_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.21 ps=1.42 w=1 l=0.15
X344 _078_ counter\[10\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X345 a_5307_4943# a_4443_4949# a_5050_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X346 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X347 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X348 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X349 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X350 VGND a_3267_9019# a_3225_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X351 a_8504_9673# a_8105_9301# a_8378_9295# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X352 a_4781_9673# a_4227_9513# a_4434_9572# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X353 VPWR a_4801_10973# a_4901_11191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X354 a_7239_8207# a_6375_8213# a_6982_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X355 _074_ a_2143_7232# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X356 _061_ a_4135_4373# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X357 a_3241_4399# a_2971_4399# a_3137_4765# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X358 VPWR net6 a_10239_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X359 a_3943_9527# a_4234_9417# a_4185_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X360 VGND counter\[3\] _050_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X361 VPWR _081_ a_5537_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X362 VGND a_7263_7637# _086_ VGND sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.10725 ps=0.98 w=0.65 l=0.15
X363 VPWR a_3593_8181# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X364 VPWR a_3819_4917# a_3735_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X365 VPWR _040_ a_5871_9527# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X366 VGND a_3593_8181# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X367 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X368 VPWR _069_ a_9965_11177# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X370 a_7607_4765# a_6909_4399# a_7350_4511# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X371 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X372 a_7102_6575# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X373 a_10103_9991# _053_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X374 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X375 VPWR a_6060_6549# _041_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X376 VGND a_6154_8863# a_6112_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X377 VGND counter\[1\] a_8205_8527# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X378 _038_ a_2509_4663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X379 a_8569_6031# _021_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X380 a_3847_9527# a_3943_9527# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X381 a_7531_2741# net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X382 VPWR net3 a_8123_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X383 VGND _031_ a_4120_3291# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10785 ps=1.36 w=0.42 l=0.15
X384 a_8102_4943# a_7663_4949# a_8017_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X385 a_2509_4663# _024_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X386 VPWR net13 _043_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X387 a_6219_4765# a_5437_4399# a_6135_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X388 a_1761_2999# net9 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X390 a_3099_9117# a_2235_8751# a_2842_8863# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X391 VGND _031_ a_7729_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X392 VGND a_4831_7093# a_4789_7497# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X393 VPWR a_5475_4917# a_5391_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X394 a_7638_7663# net3 a_7542_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X395 clknet_0_clk a_5433_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X396 a_2769_8029# a_2235_7663# a_2674_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X397 a_8397_2767# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X398 a_4009_6575# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X399 VPWR a_7407_8181# a_7323_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X400 a_5607_10089# counter\[3\] a_5513_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X401 a_6112_8751# a_5713_8751# a_5986_9117# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X402 VPWR a_6411_9117# a_6579_9019# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X403 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X404 VPWR a_9926_8181# _083_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15575 pd=1.355 as=0.135 ps=1.27 w=1 l=0.15
X405 a_8228_5321# a_7829_4949# a_8102_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X406 a_8302_7485# a_7987_7351# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X407 VGND a_3479_10004# _003_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X408 VGND a_4663_9117# a_4831_9019# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X409 _039_ net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X411 a_3593_8181# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X412 a_8017_4943# _002_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X414 VPWR _024_ a_3847_3463# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.074375 ps=0.815 w=0.42 l=0.15
X415 a_4882_4943# a_4443_4949# a_4797_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X416 VGND a_9739_6005# _036_ VGND sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X418 VPWR net10 _039_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X419 VPWR a_2439_10107# a_2355_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X420 _030_ a_4901_11191# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X421 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X422 VPWR net11 a_9777_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X423 VPWR a_7102_6575# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X424 a_5433_7637# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X425 a_2924_6575# _039_ a_2824_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X426 a_7987_7828# _077_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X427 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X428 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X429 a_9411_7119# _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X430 VGND a_2271_10205# a_2439_10107# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X431 a_8399_5487# net5 a_8293_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X432 VPWR net11 a_3042_6825# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X433 _002_ a_6375_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X434 VPWR a_3267_9019# a_3183_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X435 a_5008_5321# a_4609_4949# a_4882_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X437 a_7005_6031# _014_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X438 a_8091_10615# net8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X439 a_2229_5263# counter\[8\] a_2133_5263# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X440 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X441 VPWR a_10199_3285# net1 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X442 VPWR net10 a_6189_6825# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X443 VGND clknet_0_clk a_3593_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X444 a_4363_9673# a_4234_9417# a_3943_9527# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X445 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X446 VGND a_10199_2197# net2 VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X447 clknet_1_1__leaf_clk a_7102_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X448 counter\[0\] a_4831_7931# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X449 VPWR a_3593_8181# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X450 VPWR a_4663_9117# a_4831_9019# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X452 VGND a_7350_4511# a_7308_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X453 a_4609_4949# a_4443_4949# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X454 a_7182_4765# a_6743_4399# a_7097_4399# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X455 VPWR net7 a_9411_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X456 VPWR a_5433_7637# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X457 _026_ net7 a_5356_9615# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.091 ps=0.93 w=0.65 l=0.15
X458 _052_ net2 a_9411_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.18 ps=1.36 w=1 l=0.15
X459 a_2295_5461# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X460 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X461 clknet_0_clk a_5433_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X462 VPWR counter\[3\] a_4135_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X463 a_8727_8181# _053_ a_9158_8527# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X464 a_7641_6409# a_6651_6037# a_7515_6031# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X465 VGND _010_ a_2849_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X466 a_3226_4943# a_2953_4949# a_3141_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X467 VGND counter\[1\] _050_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X468 VPWR a_9079_6031# a_9247_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X469 VPWR _009_ a_4781_9673# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X470 a_7308_4399# a_6909_4399# a_7182_4765# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X472 counter\[0\] a_4831_7931# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X473 a_1846_10205# a_1573_9839# a_1761_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X474 _079_ a_2409_5263# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.160875 ps=1.145 w=0.65 l=0.15
X475 net12 a_2439_10107# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X476 a_3997_3317# _032_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.122275 ps=1.08 w=0.42 l=0.15
X477 _021_ a_2787_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.203125 ps=1.275 w=0.65 l=0.15
X478 _056_ counter\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X479 a_3300_9269# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X480 clknet_1_0__leaf_clk a_3593_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X481 VPWR a_6154_8863# a_6081_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X482 clknet_1_0__leaf_clk a_3593_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X483 a_4901_11191# _029_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X484 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X485 a_9739_6005# net8 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X486 VGND a_8803_9295# a_8971_9269# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X487 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X488 VGND counter\[2\] a_5633_10703# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X489 _039_ net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X490 VPWR counter\[7\] a_1559_2473# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X491 VPWR clknet_0_clk a_7102_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X492 VPWR _069_ a_3513_6825# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X493 ones[2] a_10239_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X494 a_3608_4215# a_3421_3855# a_3521_3971# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X496 VPWR a_5043_4564# _015_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X497 a_5713_8751# a_5547_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X498 a_7097_4399# _005_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X499 a_6081_9117# a_5547_8751# a_5986_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X500 clknet_1_1__leaf_clk a_7102_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X501 VGND clknet_1_1__leaf_clk a_6743_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X502 VPWR a_7625_5461# _066_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X503 VGND net7 a_9411_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X504 counter\[4\] a_3267_7931# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X505 a_5437_4399# a_5271_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X506 a_7258_6005# a_7090_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X507 VPWR a_4526_9813# a_4455_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X508 VGND _046_ a_2941_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.117 ps=1.01 w=0.65 l=0.15
X509 a_4622_6575# a_4307_6727# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X510 a_5433_7637# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X511 VPWR net11 a_9687_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X512 a_6033_9661# _041_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X513 a_8091_10615# net9 a_8265_10721# VGND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X514 a_9735_5639# net5 a_9975_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X515 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X516 VPWR a_3394_4917# a_3321_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X517 a_8574_7396# a_8367_7337# a_8750_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X518 a_2651_5487# a_2431_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X519 a_4319_9813# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X520 a_2409_5263# counter\[10\] a_2051_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X521 a_4403_6549# a_4694_6849# a_4645_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X522 a_5496_9269# _024_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X523 a_6060_6549# net11 a_6283_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X524 a_4663_8029# a_3965_7663# a_4406_7775# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X525 a_7102_6575# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X526 VGND _007_ a_4873_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X527 VPWR _057_ a_1775_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X528 a_7197_10927# _071_ a_6979_10901# VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X529 a_4047_6397# _034_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196275 ps=1.33 w=0.42 l=0.15
X530 a_4249_6397# net7 a_4143_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X531 a_3321_4943# a_2787_4949# a_3226_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X532 VPWR a_7515_6031# a_7683_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X533 a_8750_7119# a_8503_7497# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X534 _012_ _084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X535 counter\[4\] a_3267_7931# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X536 VGND a_3819_4917# a_3777_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X537 a_9975_5487# net3 a_9868_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.125125 ps=1.035 w=0.65 l=0.15
X538 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X539 clknet_1_1__leaf_clk a_7102_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X540 a_4135_4373# counter\[0\] a_4616_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X541 VGND a_3847_3463# _033_ VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X542 a_10199_3285# pulse VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X543 a_9411_7119# _051_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X544 a_9785_9661# net7 a_9713_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X545 a_9011_3285# _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.27995 ps=1.615 w=0.42 l=0.15
X546 a_5537_10703# counter\[0\] _058_ VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X547 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X548 a_2953_4949# a_2787_4949# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X549 clknet_0_clk a_5433_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X550 VGND clknet_1_1__leaf_clk a_7663_4949# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X551 a_8749_6031# a_8215_6037# a_8654_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X552 VGND counter\[2\] _050_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X553 a_6184_9839# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X554 VGND _036_ a_4981_6263# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X555 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X557 a_7749_2767# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X559 a_4406_7093# a_4238_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X560 VGND _059_ a_2665_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X561 VPWR counter\[0\] a_5607_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X562 a_9558_7775# a_9390_8029# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X563 clknet_1_0__leaf_clk a_3593_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X564 VPWR a_2271_10205# a_2439_10107# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X565 a_6729_8207# _008_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X566 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X567 a_6817_6037# a_6651_6037# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X568 VGND _053_ a_6835_5853# VGND sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.1113 ps=1.37 w=0.42 l=0.15
X569 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X570 a_4153_7663# _000_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X571 VGND net1 _081_ VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X572 _076_ _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X573 a_4675_9839# a_4455_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X574 _011_ _082_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X575 a_4415_3087# net3 a_4225_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X576 a_7917_3087# net12 a_7833_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X577 VGND net2 a_9735_5639# VGND sky130_fd_pr__nfet_01v8 ad=0.134875 pd=1.065 as=0.105625 ps=0.975 w=0.65 l=0.15
X578 a_4601_5737# counter\[3\] a_4351_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X579 a_8083_7351# a_8374_7241# a_8325_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X580 VPWR a_7102_6575# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X581 VGND net13 a_9648_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X582 VPWR a_9551_9527# _027_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X583 VPWR _024_ a_4901_11191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X584 VPWR _086_ a_5271_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X585 clknet_1_1__leaf_clk a_7102_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X586 a_10045_4943# counter\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X587 a_2502_5461# a_2302_5761# a_2651_5487# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X588 a_3353_7479# counter\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.122275 ps=1.08 w=0.42 l=0.15
X589 VGND a_6335_5461# _054_ VGND sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X590 a_5878_4511# a_5710_4765# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X591 net3 a_3819_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X592 a_8929_9673# a_7939_9301# a_8803_9295# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X594 _018_ a_2734_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X595 a_3413_4399# _050_ a_3313_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0735 ps=0.77 w=0.42 l=0.15
X596 a_6909_4399# a_6743_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X597 a_9815_8029# a_9117_7663# a_9558_7775# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X598 a_9861_5737# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1425 ps=1.285 w=1 l=0.15
X599 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X600 a_8491_3087# net3 a_8397_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X601 a_2502_5461# a_2295_5461# a_2678_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X602 VPWR counter\[0\] a_5018_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X603 VGND counter\[8\] a_10134_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X604 a_6261_4399# a_5271_4399# a_6135_4765# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X605 VPWR a_7987_7351# net6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X606 VGND clknet_0_clk a_3593_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X608 a_1751_2223# counter\[8\] a_1655_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X609 VGND _040_ a_2941_6351# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.118625 ps=1.015 w=0.65 l=0.15
X610 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X611 VPWR counter\[1\] a_8953_2473# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X612 a_9117_7663# a_8951_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X613 a_2409_5263# counter\[7\] a_2325_5263# VGND sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.08775 ps=0.92 w=0.65 l=0.15
X614 a_4663_7119# a_3965_7125# a_4406_7093# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X615 VGND a_3593_8181# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X616 VGND a_4406_7775# a_4364_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X617 a_1573_9839# a_1407_9839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X618 VGND a_9079_6031# a_9247_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X619 VGND a_9247_6005# a_9205_6409# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X620 net13 a_9983_7931# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X621 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X622 a_4238_8029# a_3799_7663# a_4153_7663# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X623 a_4153_7119# _015_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X624 a_4227_9513# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X625 a_8367_7337# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X626 a_4797_4943# _006_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X627 a_8293_9295# _022_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X628 VGND a_7711_3463# _051_ VGND sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X629 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X631 VPWR a_10103_9991# _077_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X632 VGND a_7102_6575# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X633 VGND net11 a_9687_4943# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X634 a_6154_8863# a_5986_9117# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X635 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X636 VGND a_9558_6687# a_9516_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X637 VPWR a_5871_9527# _042_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X638 a_9390_6941# a_8951_6575# a_9305_6575# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X639 a_4526_9813# a_4326_10113# a_4675_9839# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X640 net2 a_10199_2197# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X641 a_6982_8181# a_6814_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X642 VPWR clknet_1_1__leaf_clk a_6651_6037# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X643 a_3847_6727# _061_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X644 a_1761_9839# _019_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X645 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X646 a_4364_7663# a_3965_7663# a_4238_8029# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X647 a_10136_4943# _053_ a_9963_5263# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X648 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X649 clknet_1_0__leaf_clk a_3593_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X650 a_5799_9839# counter\[1\] a_5703_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X651 VPWR counter\[9\] a_2051_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X652 _059_ a_9122_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X653 clknet_1_0__leaf_clk a_3593_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X654 net13 a_9983_7931# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X655 ones[1] a_9503_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X656 a_5241_6575# a_4694_6849# a_4894_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X657 a_8653_5321# a_7663_4949# a_8527_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X658 VPWR a_3851_6005# _035_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X659 VGND a_4307_6727# net10 VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X660 a_2401_8751# a_2235_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X662 a_2011_5461# a_2302_5761# a_2253_5853# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X664 ones[10] a_9963_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X665 a_9516_6575# a_9117_6575# a_9390_6941# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X666 VGND a_3203_7351# _049_ VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X667 a_4873_9839# a_4319_9813# a_4526_9813# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X668 VGND _069_ a_1751_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X669 VGND a_6982_8181# a_6940_8585# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X670 VPWR counter\[2\] a_5607_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X671 a_4153_7663# _000_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X672 clknet_1_1__leaf_clk a_7102_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X673 VGND net14 _024_ VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X674 a_3965_7663# a_3799_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X675 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X676 a_2589_8751# _003_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X677 a_2409_4445# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X678 ones[5] a_10239_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X679 VPWR clknet_1_0__leaf_clk a_3799_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X680 VGND clknet_1_0__leaf_clk a_3799_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X681 VPWR counter\[7\] _073_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X682 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X683 a_3137_4765# a_2971_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.0567 ps=0.69 w=0.42 l=0.15
X684 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X685 a_5710_4765# a_5437_4399# a_5625_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X686 _040_ _031_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X687 VGND clk a_5433_7637# VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X688 VPWR a_8268_2741# _023_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X689 clknet_0_clk a_5433_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X690 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X691 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X692 a_3394_4917# a_3226_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X693 VPWR net6 a_8123_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X694 VPWR _083_ a_9739_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X695 VGND a_7515_6031# a_7683_6005# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X696 a_8723_7485# a_8503_7497# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X697 _068_ a_8767_10749# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X698 a_2674_8029# a_2235_7663# a_2589_7663# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X699 a_9305_6575# _018_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X700 a_4687_6549# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X701 VGND a_5433_7637# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X702 _075_ a_1465_2473# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X703 VPWR a_2295_5461# a_2302_5761# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X704 ready a_9963_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X705 a_8083_7351# a_8367_7337# a_8302_7485# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X706 a_7599_6031# a_6817_6037# a_7515_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X707 VGND a_8727_8181# _010_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X708 a_5363_6031# net3 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1475 ps=1.295 w=1 l=0.15
X709 _004_ counter\[4\] a_6184_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.091 ps=0.93 w=0.65 l=0.15
X710 VGND a_4227_9513# a_4234_9417# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X711 a_9648_2741# net12 a_9871_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X712 a_10031_6397# _083_ a_9935_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X713 VGND a_4981_6263# _037_ VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X714 a_10103_9991# _053_ a_10337_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X715 counter\[2\] a_8695_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X716 a_4238_8029# a_3965_7663# a_4153_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X718 a_9899_6941# a_9117_6575# a_9815_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X719 a_3965_7125# a_3799_7125# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X720 a_8397_2767# _083_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X721 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X722 VPWR a_3593_8181# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X723 _060_ a_2511_2223# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X724 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X725 VGND a_7102_6575# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X726 a_2014_9951# a_1846_10205# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X727 a_2431_5487# a_2302_5761# a_2011_5461# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X728 a_2800_7663# a_2401_7663# a_2674_8029# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X729 a_5050_4917# a_4882_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X730 clknet_1_1__leaf_clk a_7102_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X731 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X732 VPWR a_5433_7637# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X733 VPWR a_4894_6549# a_4823_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X734 VPWR a_5503_11092# _017_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X735 a_4238_7119# a_3799_7125# a_4153_7119# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X736 clknet_1_0__leaf_clk a_3593_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X737 a_6982_8181# a_6814_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X738 a_5271_9295# net7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X739 a_1924_2883# net9 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X740 VGND _054_ a_2879_8207# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X741 VGND a_3867_9813# counter\[7\] VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X742 a_5050_4917# a_4882_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X743 a_3099_8029# a_2401_7663# a_2842_7775# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X744 VGND clknet_1_1__leaf_clk a_6375_8213# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X745 ones[5] a_10239_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X746 VGND counter\[1\] a_7833_8903# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X747 VGND a_2842_8863# a_2800_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X748 a_2573_3087# _044_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.1365 ps=1.07 w=0.65 l=0.15
X749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X750 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X751 a_5633_10703# counter\[1\] a_5537_10703# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X752 VPWR net11 _039_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X753 a_8611_4943# a_7829_4949# a_8527_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X754 VGND _069_ a_7192_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X755 VPWR a_6579_9019# a_6495_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X756 a_1407_4399# _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X757 VPWR a_4663_7119# a_4831_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X759 a_4364_7497# a_3965_7125# a_4238_7119# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X760 a_9926_8181# net14 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10675 ps=1.005 w=0.42 l=0.15
X761 VGND a_9011_3285# _031_ VGND sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.10725 ps=0.98 w=0.65 l=0.15
X762 VPWR a_5307_4943# a_5475_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X763 a_4747_9117# a_3965_8751# a_4663_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X764 counter\[5\] a_7775_4667# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X765 a_3421_3855# _065_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X766 a_3651_4943# a_2787_4949# a_3394_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X767 VPWR a_4406_7775# a_4333_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X768 a_7733_4399# a_6743_4399# a_7607_4765# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X769 a_4589_3829# net8 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X770 a_3593_8181# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X771 VGND a_7775_4667# a_7733_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X772 VPWR a_8803_9295# a_8971_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X773 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X775 a_4687_6549# clknet_1_1__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X776 VPWR a_7239_8207# a_7407_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X778 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X779 a_4238_7119# a_3965_7125# a_4153_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X780 a_3434_7479# counter\[10\] a_3353_7479# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.05355 ps=0.675 w=0.42 l=0.15
X781 VPWR clknet_1_1__leaf_clk a_8951_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X782 a_10048_10927# _069_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X783 _064_ a_10136_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X784 a_9899_8029# a_9117_7663# a_9815_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X785 a_4333_8029# a_3799_7663# a_4238_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X786 a_2674_8029# a_2401_7663# a_2589_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X787 VGND _069_ a_6093_8527# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X788 a_10141_8323# net14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.15575 ps=1.355 w=0.42 l=0.15
X789 VPWR _007_ a_4873_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X790 VPWR net9 a_8091_10615# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X791 VGND a_9983_6843# a_9941_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X792 clknet_0_clk a_5433_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X793 a_8378_9295# a_8105_9301# a_8293_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X794 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X795 VPWR a_7531_2741# _047_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X796 a_4455_9839# a_4326_10113# a_4035_9813# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X797 VGND a_5503_11092# _017_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X798 a_9739_6005# net9 a_10137_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X799 a_9043_10749# counter\[6\] a_8937_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X800 VGND a_6411_9117# a_6579_9019# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X801 a_2589_8751# _003_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X802 a_8205_5487# net7 a_8123_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X803 a_6979_10901# _071_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X804 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X805 _005_ a_5823_7119# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X806 a_7263_7637# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07455 pd=0.775 as=0.0777 ps=0.79 w=0.42 l=0.15
X807 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X808 _028_ a_8123_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X809 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X810 VPWR clknet_1_1__leaf_clk a_8951_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X811 _044_ net12 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X812 _008_ a_5731_3311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X813 VGND _013_ a_8921_7497# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X815 VPWR a_4589_3829# _029_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X816 a_9551_9527# net8 a_9785_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X817 a_4601_5737# counter\[2\] a_4798_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X818 a_8197_4943# a_7663_4949# a_8102_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X819 VPWR _010_ a_2849_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X820 VGND a_8695_4917# a_8653_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X821 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X822 _050_ a_5018_5461# a_4798_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X823 a_3042_6825# _035_ a_2734_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X824 ones[8] a_9687_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X825 a_4319_2767# _080_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X826 VPWR _062_ a_7343_7351# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.074375 ps=0.815 w=0.42 l=0.15
X827 VPWR net11 a_7749_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X828 VPWR a_4406_7093# a_4333_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X829 _039_ net11 a_7479_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X830 VPWR clknet_1_1__leaf_clk a_7939_9301# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X831 VGND net2 _024_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X832 VPWR net10 a_3851_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0735 ps=0.77 w=0.42 l=0.15
X833 VPWR a_2842_7775# a_2769_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X834 _080_ net14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X835 VGND a_7102_6575# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X836 VPWR a_8546_9269# a_8473_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X837 _052_ _049_ a_9661_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.0975 ps=0.95 w=0.65 l=0.15
X838 a_7479_10927# net10 a_7729_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X839 VPWR _066_ a_3521_3971# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X840 clknet_1_0__leaf_clk a_3593_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X841 VPWR a_2439_10107# net12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X842 a_7928_5487# counter\[4\] a_7625_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X843 VPWR a_7102_6575# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X844 a_2133_5263# _069_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X845 VPWR a_5433_7637# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X846 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X847 a_9935_6397# _028_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.196275 ps=1.33 w=0.42 l=0.15
X848 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X849 a_4333_7119# a_3799_7125# a_4238_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X850 a_7097_4399# _005_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X851 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X852 a_6335_5461# a_6511_5461# a_6463_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X853 VPWR a_8355_4074# _022_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X854 a_4977_4943# a_4443_4949# a_4882_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X855 a_2824_6575# _024_ a_2734_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X856 a_8473_9295# a_7939_9301# a_8378_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X857 net3 a_3819_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X858 _083_ a_9926_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X859 a_4491_6263# _056_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X860 VPWR a_1673_10973# a_1773_11191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X861 VPWR a_7607_4765# a_7775_4667# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X862 a_9205_6409# a_8215_6037# a_9079_6031# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X863 _014_ a_2776_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.3275 ps=1.655 w=1 l=0.15
X864 a_7108_5737# a_6835_5853# _071_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X865 VPWR a_7833_8903# _055_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X866 a_4801_10973# _027_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X867 VGND a_3847_9527# counter\[9\] VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X868 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X869 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X870 _026_ a_5496_9269# a_5271_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X871 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X872 a_1573_9839# a_1407_9839# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X873 clknet_1_1__leaf_clk a_7102_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X874 a_6189_6575# _036_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X875 a_7833_8903# counter\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X876 VGND clknet_1_1__leaf_clk a_8951_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X877 VPWR a_3593_8181# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X878 ones[6] a_9043_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X879 ones[8] a_9687_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X880 a_7833_8903# counter\[1\] a_7996_9001# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X881 _004_ a_6324_10029# a_6099_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X882 a_9735_5639# net14 a_10204_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=1.415 w=1 l=0.15
X883 clknet_0_clk a_5433_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X884 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X885 VPWR net1 a_4319_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X886 VGND a_10103_9991# _077_ VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X887 a_9011_3285# net9 a_9492_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06195 ps=0.715 w=0.42 l=0.15
X888 VPWR a_2502_5461# a_2431_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X889 VGND a_5433_7637# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X890 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X891 a_2953_4949# a_2787_4949# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X892 _053_ a_3300_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X893 VGND a_7607_4765# a_7775_4667# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X894 VPWR a_6612_3829# _069_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X895 a_8727_8181# _076_ a_8945_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X896 a_2769_9117# a_2235_8751# a_2674_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X897 VGND net13 _043_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X898 a_1559_2473# counter\[9\] a_1465_2473# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X899 VPWR counter\[0\] a_4135_4373# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07455 ps=0.775 w=0.42 l=0.15
X900 ones[2] a_10239_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X902 a_9661_7439# _050_ a_9411_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X903 _076_ counter\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X904 VGND a_4135_4373# _061_ VGND sky130_fd_pr__nfet_01v8 ad=0.17515 pd=1.265 as=0.10725 ps=0.98 w=0.65 l=0.15
X905 a_9117_4399# net10 a_9033_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X906 a_8075_3285# counter\[7\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X907 VPWR clknet_1_0__leaf_clk a_2235_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X908 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X909 VGND clknet_1_0__leaf_clk a_2235_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X910 a_5307_4943# a_4609_4949# a_5050_4917# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X911 a_8105_9301# a_7939_9301# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X912 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X913 _082_ a_4225_2767# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X914 VPWR a_7987_7828# _009_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X915 a_7749_2767# net4 a_7531_2741# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X916 _073_ counter\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X917 a_9158_8527# _079_ a_8863_8527# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X918 a_5529_7439# counter\[8\] a_5445_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X919 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X920 VGND a_4663_7119# a_4831_7093# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X921 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X922 VPWR counter\[10\] a_3203_7351# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.074375 ps=0.815 w=0.42 l=0.15
X923 VPWR _073_ a_2143_7232# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X924 _070_ _065_ a_1489_4649# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X925 VGND net7 a_2603_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X926 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X927 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X928 VGND a_7239_8207# a_7407_8181# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X929 VPWR net4 _046_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X930 a_3183_8029# a_2401_7663# a_3099_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X931 a_7729_10927# net10 a_7479_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X932 VPWR a_9735_5639# _085_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.285 ps=2.57 w=1 l=0.15
X933 a_4789_7663# a_3799_7663# a_4663_8029# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X934 VGND _017_ a_5241_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X935 VPWR net14 a_8231_4649# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X936 _067_ a_3521_3971# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X937 a_5871_9527# _024_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X938 _046_ net4 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X939 VPWR _031_ a_4120_3291# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1087 ps=1.36 w=0.42 l=0.15
X940 VGND a_4831_7931# a_4789_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X941 a_9558_6687# a_9390_6941# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X942 a_9551_9527# _086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X943 _008_ a_5731_3311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X944 a_7711_3463# counter\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X945 a_3137_4765# _050_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1281 ps=1.03 w=0.42 l=0.15
X946 a_7493_7479# _052_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.122275 ps=1.08 w=0.42 l=0.15
X947 VGND a_10199_3285# net1 VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X948 VGND a_8270_4917# a_8228_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X949 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X950 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X951 _078_ counter\[10\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X952 VPWR clknet_1_0__leaf_clk a_1407_9839# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X953 VPWR _060_ a_6375_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X954 a_3203_7351# counter\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.142225 ps=1.335 w=0.42 l=0.15
X955 a_8654_6031# a_8381_6037# a_8569_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X956 a_4873_9839# a_4326_10113# a_4526_9813# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X957 a_9941_6575# a_8951_6575# a_9815_6941# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X958 VPWR _061_ a_6099_10089# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X959 VPWR a_2007_7828# _019_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X960 VPWR clknet_0_clk a_3593_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X961 VGND _027_ a_1761_2999# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X962 a_4707_10703# net3 _084_ VGND sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X963 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X964 a_9965_11177# counter\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X965 a_8381_6037# a_8215_6037# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X966 a_2842_7775# a_2674_8029# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X967 a_6612_3829# _068_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X968 a_4225_2767# net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X969 VGND _061_ a_7928_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X970 a_6060_6549# net12 a_6189_6825# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X971 a_7691_4765# a_6909_4399# a_7607_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X972 a_5043_6575# a_4823_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X973 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X974 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X975 net5 a_4831_9019# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X976 VPWR a_5433_7637# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X977 a_3847_3463# a_4120_3291# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1085 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X978 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X979 a_1761_2999# _027_ a_1924_2883# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X980 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X981 VPWR _067_ a_5823_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X982 VPWR a_4434_9572# a_4363_9673# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X983 a_2271_10205# a_1407_9839# a_2014_9951# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X984 VPWR counter\[7\] a_7108_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X985 VPWR net12 _044_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X986 VPWR counter\[7\] a_7282_11177# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X987 ones[9] a_9687_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X988 _040_ net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X989 _069_ a_6612_3829# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X990 VPWR a_8822_6005# a_8749_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X991 VGND a_5307_4943# a_5475_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X992 VGND a_7102_6575# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X993 a_3479_10004# _063_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X994 a_5713_8751# a_5547_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X995 a_5871_9527# _041_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.142225 ps=1.335 w=0.42 l=0.15
X996 net12 a_2439_10107# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X997 ones[6] a_9043_5487# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X998 a_9963_5263# _061_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X999 VPWR a_7683_6005# net7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1000 a_4653_6397# _056_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X1001 clknet_1_0__leaf_clk a_3593_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1002 a_1655_2223# counter\[7\] a_1465_2473# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1003 VPWR a_5433_7637# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1004 VPWR a_2014_9951# a_1941_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1005 VPWR a_3847_6727# _065_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X1006 VGND a_9648_2741# _045_ VGND sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1007 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1008 a_4823_6575# a_4694_6849# a_4403_6549# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1009 a_4789_7497# a_3799_7125# a_4663_7119# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1010 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1011 VGND _051_ a_9411_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1012 VGND a_7343_7351# _063_ VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.169 ps=1.82 w=0.65 l=0.15
X1013 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1015 VGND a_5018_5461# _050_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1016 VPWR a_3867_9813# counter\[7\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1017 a_4797_4943# _006_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1018 a_4663_9117# a_3965_8751# a_4406_8863# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1019 VPWR a_4831_7931# counter\[0\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1020 VGND _061_ a_7616_7351# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10785 ps=1.36 w=0.42 l=0.15
X1021 VGND _028_ a_4892_4175# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1022 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1023 VPWR clknet_1_1__leaf_clk a_8215_6037# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1024 VGND a_8822_6005# a_8780_6409# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1025 a_9305_6575# _018_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1026 VGND a_7987_7828# _009_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1027 a_4621_10383# net5 _084_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1028 VGND a_5878_4511# a_5836_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1029 a_7277_4765# a_6743_4399# a_7182_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1030 net5 a_4831_9019# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1031 a_3313_4399# _049_ a_3241_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0441 ps=0.63 w=0.42 l=0.15
X1032 a_5710_4765# a_5271_4399# a_5625_4399# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1033 a_9777_3087# _035_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1034 a_3847_6727# counter\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1035 counter\[3\] a_3267_9019# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1036 clknet_0_clk a_5433_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1037 a_4162_9661# a_3847_9527# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X1038 a_2501_3087# _024_ a_2419_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X1039 _062_ a_5513_10089# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X1040 ones[9] a_9687_10927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1041 a_2051_4943# counter\[8\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1042 a_4894_6549# a_4694_6849# a_5043_6575# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1043 _074_ a_2143_7232# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1044 VGND a_3593_8181# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1045 VPWR a_4307_6727# net10 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1046 a_5060_10933# _029_ a_4988_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X1047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1048 a_5878_4511# a_5710_4765# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1049 ones[10] a_9963_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1050 a_5836_4399# a_5437_4399# a_5710_4765# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1051 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1052 a_4894_6549# a_4687_6549# a_5070_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X1053 _024_ net2 a_8231_4649# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1054 a_7192_5487# counter\[7\] _071_ VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X1055 VPWR counter\[1\] _056_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1056 VGND a_8355_4074# _022_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1057 a_5241_6575# a_4687_6549# a_4894_6549# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1058 VPWR a_7407_8181# counter\[8\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1059 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1060 a_6463_5487# _053_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X1061 net14 a_8971_9269# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1063 a_4153_8751# _012_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1064 a_5070_6941# a_4823_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X1065 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1066 a_7843_5737# counter\[5\] a_7625_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1068 a_8569_6031# _021_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1069 _040_ net12 a_9201_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X1070 ready a_9963_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1071 _031_ a_9011_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X1072 a_6729_8207# _008_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1073 _052_ net2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X1074 a_6909_4399# a_6743_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1075 a_9163_6031# a_8381_6037# a_9079_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1076 a_2869_6351# _024_ a_2787_6031# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X1077 VGND a_2007_7828# _019_ VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1078 a_9305_7663# _020_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1079 VPWR _024_ a_1773_11191# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1080 VPWR clk a_5433_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1081 _079_ a_2409_5263# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1082 counter\[3\] a_3267_9019# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1083 _076_ counter\[7\] a_5613_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X1084 a_10137_6397# net8 a_10031_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.0798 ps=0.8 w=0.42 l=0.15
X1085 VPWR net9 a_9011_3285# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07455 ps=0.775 w=0.42 l=0.15
X1086 VPWR a_9739_6005# _036_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.26 ps=2.52 w=1 l=0.15
X1087 _043_ net13 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1088 a_6135_4765# a_5271_4399# a_5878_4511# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1089 clknet_1_1__leaf_clk a_7102_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1090 _016_ a_5271_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1091 VPWR _061_ a_8767_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1092 VGND net4 a_9963_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1093 a_5043_4564# _030_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1094 a_7574_7479# _062_ a_7493_7479# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.05355 ps=0.675 w=0.42 l=0.15
X1095 counter\[7\] a_3867_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1096 VGND a_5433_7637# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1097 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1098 a_8123_5487# net7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X1099 clknet_0_clk a_5433_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1100 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1101 a_8075_3285# counter\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1102 a_6541_8213# a_6375_8213# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1103 a_7263_7637# net1 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.27995 ps=1.615 w=0.42 l=0.15
X1104 a_4621_10383# _083_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X1105 VPWR _053_ a_2143_7232# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1106 net7 a_7683_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1107 VGND a_4491_6263# _057_ VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1108 VGND _085_ _012_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1109 VGND counter\[8\] a_3476_7351# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10785 ps=1.36 w=0.42 l=0.15
X1110 VGND a_4406_8863# a_4364_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1111 a_7108_5737# _069_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1112 a_4238_9117# a_3799_8751# a_4153_8751# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1113 VPWR clknet_0_clk a_3593_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1114 a_2225_7485# _053_ a_2143_7232# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1115 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1116 a_9036_2223# counter\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1117 VGND counter\[6\] a_1407_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1119 VPWR _059_ a_2511_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X1120 VGND net6 a_8268_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1121 VPWR a_3593_8181# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1122 _001_ a_1775_4399# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1123 a_7005_6031# _014_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1124 VGND clknet_0_clk a_7102_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1125 VGND a_9558_7775# a_9516_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1126 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1127 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1128 a_2776_7119# _026_ a_2603_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1129 a_9390_8029# a_8951_7663# a_9305_7663# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1130 VPWR a_6303_4667# a_6219_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1131 net1 a_10199_3285# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1132 a_4364_8751# a_3965_8751# a_4238_9117# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1133 a_1846_10205# a_1407_9839# a_1761_9839# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1134 VGND a_7683_6005# net7 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1135 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1136 a_3394_4917# a_3226_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1137 VPWR a_8367_7337# a_8374_7241# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1138 a_6411_9117# a_5547_8751# a_6154_8863# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1139 _016_ a_5271_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1140 net2 a_10199_2197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1141 a_7479_10927# net11 _039_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1143 VGND _043_ a_2573_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.117 ps=1.01 w=0.65 l=0.15
X1144 a_4351_5737# counter\[3\] a_4601_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1145 VPWR a_7263_7637# _086_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.165 ps=1.33 w=1 l=0.15
X1146 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1147 VPWR a_9983_6843# net11 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1148 VGND counter\[2\] a_5799_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X1149 a_9516_7663# a_9117_7663# a_9390_8029# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1150 a_6154_8863# a_5986_9117# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1151 a_3867_9813# a_4035_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1152 a_8727_8181# _053_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X1153 _006_ _070_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1154 clknet_1_0__leaf_clk a_3593_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1155 a_4153_8751# _012_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1156 a_1972_9839# a_1573_9839# a_1846_10205# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1157 _048_ a_3137_4765# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1034 ps=1 w=0.65 l=0.15
X1158 VGND _060_ a_6375_2767# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1159 a_7350_4511# a_7182_4765# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1160 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1161 _086_ a_7263_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X1162 VGND clknet_1_0__leaf_clk a_3799_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1163 VGND a_2295_5461# a_2302_5761# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1164 _021_ a_2787_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3125 ps=1.625 w=1 l=0.15
X1165 _038_ a_2509_4663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1166 a_1941_10205# a_1407_9839# a_1846_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1167 a_1773_11191# _023_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X1168 a_2674_9117# a_2235_8751# a_2589_8751# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1169 _062_ a_5513_10089# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X1170 a_9305_7663# _020_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1171 a_6814_8207# a_6375_8213# a_6729_8207# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1172 a_8102_4943# a_7829_4949# a_8017_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1173 a_5607_10089# counter\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X1174 VPWR clknet_1_1__leaf_clk a_5271_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1175 VPWR net3 a_4319_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1176 a_7749_2767# net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X1177 a_1761_9839# _019_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1178 VPWR a_7258_6005# a_7185_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1179 a_9648_2741# net13 a_9777_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1180 VPWR counter\[4\] a_8767_10749# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1181 VGND a_9983_6843# net11 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1182 a_8953_2473# counter\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1183 a_3680_4215# _053_ a_3608_4215# VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X1184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1185 a_5446_6351# _080_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.17225 ps=1.83 w=0.65 l=0.15
X1186 clknet_0_clk a_5433_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1187 a_4238_9117# a_3965_8751# a_4153_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1188 _050_ counter\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1189 VPWR a_9558_6687# a_9485_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1190 VPWR _026_ a_2776_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.195 ps=1.39 w=1 l=0.15
X1191 a_6105_9661# _040_ a_6033_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1192 a_7933_3311# counter\[5\] a_7845_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X1193 VPWR _046_ a_3158_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.18 ps=1.36 w=1 l=0.15
X1194 VGND a_9551_9527# _027_ VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1195 a_6940_8585# a_6541_8213# a_6814_8207# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1196 a_2800_8751# a_2401_8751# a_2674_9117# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1198 a_7185_6031# a_6651_6037# a_7090_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1199 VPWR clknet_1_0__leaf_clk a_5547_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1200 VGND _024_ a_5060_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X1201 a_8937_10749# counter\[4\] a_8849_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1202 VGND a_7407_8181# counter\[8\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1203 _060_ a_2511_2223# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X1204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1205 a_7542_7663# net1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.17515 ps=1.265 w=0.42 l=0.15
X1206 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1207 VPWR net3 a_8397_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1208 ones[1] a_9503_8207# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1209 VGND net14 _080_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1210 a_7744_7663# net5 a_7638_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0798 ps=0.8 w=0.42 l=0.15
X1211 VPWR a_3099_8029# a_3267_7931# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1212 a_9485_6941# a_8951_6575# a_9390_6941# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1213 a_4882_4943# a_4609_4949# a_4797_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1214 VPWR clknet_1_0__leaf_clk a_3799_7125# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1215 a_3099_9117# a_2401_8751# a_2842_8863# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1216 a_7239_8207# a_6541_8213# a_6982_8181# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1217 a_5433_7637# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1218 a_2734_6575# _039_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X1219 a_9386_3311# net7 a_9290_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X1220 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1221 VGND net8 a_10239_10383# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1222 ones[4] a_10239_10383# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1223 VPWR a_8270_4917# a_8197_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1224 a_2051_4943# counter\[7\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1225 a_3851_6005# net7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0777 ps=0.79 w=0.42 l=0.15
X1226 clknet_1_0__leaf_clk a_3593_8181# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1227 VPWR net3 a_7263_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X1228 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1229 a_4078_3317# _024_ a_3997_3317# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.05355 ps=0.675 w=0.42 l=0.15
X1230 VGND a_7102_6575# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1231 a_7282_11177# _069_ a_6979_10901# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X1232 VGND net3 a_9779_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1233 VPWR a_4406_8863# a_4333_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1234 VPWR _017_ a_5241_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X1235 VGND a_3099_8029# a_3267_7931# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1237 a_7829_4949# a_7663_4949# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1238 a_2776_7119# _086_ a_2685_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1525 ps=1.305 w=1 l=0.15
X1239 VPWR a_6511_5461# a_6335_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1240 a_3965_8751# a_3799_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1241 a_3965_7663# a_3799_7663# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1242 a_4277_10205# a_3867_9813# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X1243 VPWR a_3300_9269# _053_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1244 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1245 a_3593_8181# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1246 a_4333_9117# a_3799_8751# a_4238_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1247 _061_ a_4135_4373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X1248 VPWR a_9558_7775# a_9485_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1249 VGND _078_ a_8863_8527# VGND sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1250 a_2674_9117# a_2401_8751# a_2589_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1251 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1252 VGND _039_ a_2573_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.118625 ps=1.015 w=0.65 l=0.15
X1253 VGND a_9983_7931# a_9941_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1254 VPWR clknet_1_0__leaf_clk a_2787_4949# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1255 net7 a_7683_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1256 VGND a_5871_9527# _042_ VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.169 ps=1.82 w=0.65 l=0.15
X1257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1258 _081_ net1 a_5363_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1259 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1260 a_6909_8207# a_6375_8213# a_6814_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1261 a_7102_6575# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1262 net9 a_6303_4667# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1263 _020_ a_2419_2767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.203125 ps=1.275 w=0.65 l=0.15
X1264 VGND a_6060_6549# _041_ VGND sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1265 a_4227_9513# clknet_1_0__leaf_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1266 a_9485_8029# a_8951_7663# a_9390_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1267 a_2573_3087# _045_ a_2501_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.06825 ps=0.86 w=0.65 l=0.15
X1268 a_7343_7351# _052_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.142225 ps=1.335 w=0.42 l=0.15
X1269 clknet_0_clk a_5433_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1270 a_5433_5321# a_4443_4949# a_5307_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1271 a_4981_6263# net10 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1272 VGND _009_ a_4781_9673# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X1273 a_10199_2197# rst VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1274 a_4351_5737# counter\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1276 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1277 VGND clknet_1_1__leaf_clk a_6651_6037# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1278 VPWR a_9815_6941# a_9983_6843# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1279 _000_ a_2879_8207# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1280 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1281 VPWR clknet_1_0__leaf_clk a_4443_4949# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1282 VGND a_3593_8181# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1283 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1284 a_3651_4943# a_2953_4949# a_3394_4917# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1285 VPWR _013_ a_8921_7497# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X1286 a_7833_3087# net13 a_7531_2741# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X1287 VPWR a_2842_8863# a_2769_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1288 VPWR a_3651_4943# a_3819_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1289 a_5144_6147# net10 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X1290 net9 a_6303_4667# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1291 VPWR a_3421_3855# a_3521_3971# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X1292 a_3044_6031# _040_ a_2787_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.1375 ps=1.275 w=1 l=0.15
X1293 a_9777_2767# net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1295 VGND _024_ a_1932_10933# VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X1296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1297 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1298 VGND a_6979_10901# _007_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1299 clknet_1_1__leaf_clk a_7102_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1300 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1301 _070_ _053_ a_1407_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1302 net8 a_4831_7093# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1303 a_4185_9295# a_3847_9527# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X1304 a_2355_10205# a_1573_9839# a_2271_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1305 a_9122_2223# counter\[2\] a_8953_2473# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X1306 counter\[6\] a_5475_4917# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1307 VGND a_9815_6941# a_9983_6843# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1308 a_3735_4943# a_2953_4949# a_3651_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1309 VPWR a_4319_9813# a_4326_10113# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1311 VGND a_7102_6575# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1312 net14 a_8971_9269# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1313 a_2401_7663# a_2235_7663# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1314 a_4892_4175# _083_ a_4589_3829# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1315 a_9861_5737# net5 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.305 ps=1.61 w=1 l=0.15
X1316 a_4583_9661# a_4363_9673# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X1317 VGND clknet_1_0__leaf_clk a_1407_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1318 VPWR a_8091_10615# _034_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1319 VPWR _053_ a_2511_2223# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1320 _072_ a_10134_10927# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1321 a_2924_6575# net11 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X1322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1323 VPWR _055_ a_4491_6263# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X1324 a_3943_9527# a_4227_9513# a_4162_9661# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1325 a_2790_2767# _044_ a_2676_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.21 ps=1.42 w=1 l=0.15
X1326 a_6189_6825# net11 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1327 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1328 a_4406_7775# a_4238_8029# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1329 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1330 a_4406_7775# a_4238_8029# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1331 VGND clknet_1_1__leaf_clk a_8951_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1332 a_1673_10973# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1333 a_8767_10749# counter\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X1334 a_7343_7351# a_7616_7351# a_7574_7479# VGND sky130_fd_pr__nfet_01v8 ad=0.107825 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1335 a_4510_4399# counter\[3\] a_4414_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0693 ps=0.75 w=0.42 l=0.15
X1336 counter\[1\] a_6579_9019# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1337 VGND counter\[10\] _078_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1338 a_5391_4943# a_4609_4949# a_5307_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1339 a_6283_6575# net10 a_6189_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1340 a_3421_3855# _065_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1342 a_4807_3855# net8 a_4589_3829# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1343 clknet_1_1__leaf_clk a_7102_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1344 VPWR a_3203_7351# _049_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X1345 VPWR _049_ a_3137_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.0987 ps=0.89 w=0.42 l=0.15
X1346 a_4363_9673# a_4227_9513# a_3943_9527# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X1347 VGND _066_ a_3680_4215# VGND sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X1348 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1349 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1350 a_8033_3311# counter\[6\] a_7933_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X1351 a_7515_6031# a_6817_6037# a_7258_6005# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1352 a_2941_6351# _043_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.1365 ps=1.07 w=0.65 l=0.15
X1353 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1354 a_2297_7485# _072_ a_2225_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1355 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1356 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1357 clknet_0_clk a_5433_7637# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1358 a_10134_10927# counter\[7\] a_10048_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1359 a_4798_5737# counter\[2\] a_4601_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1360 VGND clknet_1_0__leaf_clk a_2235_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1361 a_8546_9269# a_8378_9295# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1362 a_3479_10004# _063_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1363 a_1465_2473# counter\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X1364 VGND a_5433_7637# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1365 VGND counter\[0\] a_6511_5461# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1366 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1367 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1368 VPWR a_8727_8181# _010_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1369 a_3847_3463# _032_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.142225 ps=1.335 w=0.42 l=0.15
X1370 counter\[2\] a_8695_4917# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1371 a_5537_5737# _082_ _011_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1372 VGND _061_ a_9043_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1373 a_10204_5737# net2 a_9861_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.415 as=0.1625 ps=1.325 w=1 l=0.15
X1374 VGND a_3593_8181# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1375 a_8270_4917# a_8102_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1376 VPWR a_4981_6263# _037_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X1377 VGND a_8546_9269# a_8504_9673# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1378 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1379 a_7197_10927# counter\[7\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1380 a_3183_9117# a_2401_8751# a_3099_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1381 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1382 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1383 a_3226_4943# a_2787_4949# a_3141_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1384 clknet_1_1__leaf_clk a_7102_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1385 a_4789_8751# a_3799_8751# a_4663_9117# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1386 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1387 a_2842_7775# a_2674_8029# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1388 a_8574_7396# a_8374_7241# a_8723_7485# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X1389 a_8270_4917# a_8102_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1390 VPWR net5 a_9503_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1391 VPWR a_6335_5461# _054_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X1392 a_7182_4765# a_6909_4399# a_7097_4399# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1393 counter\[1\] a_6579_9019# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1394 VGND a_6324_10029# _004_ VGND sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.143 ps=1.09 w=0.65 l=0.15
X1395 a_4406_7093# a_4238_7119# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1396 VGND clknet_0_clk a_7102_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1397 _064_ a_10136_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.3275 ps=1.655 w=1 l=0.15
X1398 a_4663_8029# a_3799_7663# a_4406_7775# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1399 VPWR a_4687_6549# a_4694_6849# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1400 _018_ a_2734_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1401 VGND a_4831_9019# a_4789_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1402 a_8546_9269# a_8378_9295# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1403 VPWR net13 a_9687_10927# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1404 a_9558_7775# a_9390_8029# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1405 VPWR a_3479_10004# _003_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1406 VGND a_7407_8181# a_7365_8585# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1408 VGND a_7625_5461# _066_ VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1409 a_3352_5321# a_2953_4949# a_3226_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1410 VPWR _049_ a_9411_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.41 pd=1.82 as=0.135 ps=1.27 w=1 l=0.15
X1411 VGND a_9926_8181# _083_ VGND sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1412 VPWR a_8527_4943# a_8695_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1413 a_8921_7497# a_8367_7337# a_8574_7396# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X1414 VPWR net7 a_9551_9527# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.06615 ps=0.735 w=0.42 l=0.15
X1415 VGND a_1761_2999# _032_ VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1416 VPWR counter\[5\] a_7711_3463# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X1417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1418 VPWR _069_ a_2051_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1419 a_5433_7637# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1420 VPWR _051_ a_3137_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.06615 ps=0.735 w=0.42 l=0.15
X1421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1422 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1423 counter\[7\] a_3867_9813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1424 a_9941_7663# a_8951_7663# a_9815_8029# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1425 a_5503_11092# _038_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1426 a_10103_9514# _025_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1427 ones[3] a_9411_8751# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1428 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1429 VGND net14 a_9963_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1430 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1431 a_8527_4943# a_7663_4949# a_8270_4917# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1432 a_7102_6575# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X1433 a_3203_7351# a_3476_7351# a_3434_7479# VGND sky130_fd_pr__nfet_01v8 ad=0.107825 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1434 a_8293_9295# _022_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1435 a_5871_9527# _024_ a_6105_9661# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1437 a_2842_8863# a_2674_9117# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1438 a_9926_8181# net1 a_10141_8323# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1439 a_5901_8751# _001_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1440 VPWR a_7350_4511# a_7277_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1441 a_9411_7439# _050_ a_9661_7439# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1442 VGND clknet_1_1__leaf_clk a_7939_9301# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1443 VPWR a_7102_6575# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1444 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1445 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1446 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1447 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1448 VPWR a_4831_7931# a_4747_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1450 VPWR _069_ _073_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1451 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1452 clknet_1_1__leaf_clk a_7102_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X1454 VGND net13 a_9687_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1455 net8 a_4831_7093# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1456 a_4663_7119# a_3799_7125# a_4406_7093# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1457 VGND a_4687_6549# a_4694_6849# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1458 VGND a_8574_7396# a_8503_7497# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X1459 VPWR net4 a_9963_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1460 a_2603_7439# _086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X1461 a_8803_9295# a_7939_9301# a_8546_9269# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1462 a_5043_4564# _030_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1463 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1464 a_5703_9839# counter\[0\] a_5513_10089# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1465 a_5503_11092# _038_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1466 VPWR a_8695_4917# a_8611_4943# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1467 ones[3] a_9411_8751# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1468 a_4801_10973# _027_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1469 VGND _069_ a_7197_10927# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X1470 clknet_1_1__leaf_clk a_7102_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1471 a_8231_4649# net14 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1472 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1473 VPWR clk a_5433_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1474 _050_ counter\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1475 net4 a_9247_6005# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1476 VGND a_7102_6575# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1477 ones[7] a_9687_4943# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1478 VGND net2 _052_ VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.117 ps=1.01 w=0.65 l=0.15
X1479 VGND a_4831_7931# counter\[0\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1480 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1481 a_4645_6941# a_4307_6727# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X1482 a_5625_4399# _016_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1483 VPWR net3 a_9861_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X1484 a_10265_9839# _076_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.13165 ps=1.14 w=0.42 l=0.15
X1485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1486 a_8268_2741# net5 a_8491_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1487 VPWR a_5433_7637# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1488 a_5986_9117# a_5547_8751# a_5901_8751# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1489 a_9411_7119# _049_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.41 ps=1.82 w=1 l=0.15
X1490 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1491 VGND net2 a_2971_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1492 a_6135_4765# a_5437_4399# a_5878_4511# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1493 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1494 a_8822_6005# a_8654_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1495 _001_ a_1775_4399# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1496 a_8205_8527# counter\[0\] _056_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1497 VPWR a_4831_7093# a_4747_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1498 VPWR a_3847_9527# counter\[9\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1499 a_3851_6005# net10 a_4249_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X1500 a_2596_4405# a_2409_4445# a_2509_4663# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X1501 VPWR a_8971_9269# a_8887_9295# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1502 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1503 VPWR a_7102_6575# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1504 VPWR a_2409_4445# a_2509_4663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X1505 a_8503_7497# a_8374_7241# a_8083_7351# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X1506 a_9871_3087# net11 a_9777_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1507 clknet_1_0__leaf_clk a_3593_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1508 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1509 VGND _067_ a_5823_7119# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1510 VGND a_2502_5461# a_2431_5487# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X1511 VGND a_7683_6005# a_7641_6409# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1512 VPWR _074_ a_5731_3311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1513 VPWR a_3593_8181# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1514 _039_ _031_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1515 a_4823_6575# a_4687_6549# a_4403_6549# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X1516 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1517 a_5901_8751# _001_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1518 VGND a_5050_4917# a_5008_5321# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1519 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1520 VPWR net12 a_9687_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1521 a_3851_6005# _034_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.31245 ps=1.68 w=0.42 l=0.15
X1522 a_6411_9117# a_5713_8751# a_6154_8863# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1523 a_1505_7119# _084_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1524 VPWR _037_ a_2509_4663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1525 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1526 a_3225_7663# a_2235_7663# a_3099_8029# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1527 a_8527_4943# a_7829_4949# a_8270_4917# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1528 VGND a_2439_10107# net12 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1529 a_7829_4949# a_7663_4949# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1530 a_4319_2767# net2 a_4225_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X1531 VGND a_3593_8181# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1532 a_2014_9951# a_1846_10205# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1533 VPWR _050_ a_9411_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1534 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1535 VGND a_3267_7931# a_3225_7663# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1536 VGND clknet_1_0__leaf_clk a_2787_4949# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1537 _031_ a_9011_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.195 ps=1.9 w=0.65 l=0.15
X1538 a_10103_9514# _025_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1539 a_7711_3463# counter\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X1540 VPWR _079_ a_8727_8181# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X1541 a_5986_9117# a_5713_8751# a_5901_8751# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1542 a_9411_7439# _051_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1543 VPWR counter\[8\] _076_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1544 VGND _051_ a_3413_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.0609 ps=0.71 w=0.42 l=0.15
X1545 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1546 a_8822_6005# a_8654_6031# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1547 VGND a_4526_9813# a_4455_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X1548 _069_ a_6612_3829# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1549 a_7090_6031# a_6817_6037# a_7005_6031# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1550 _043_ net13 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1551 a_2685_7119# net7 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X1552 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1553 VPWR a_4663_8029# a_4831_7931# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1554 VPWR counter\[2\] _058_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1555 VPWR net8 a_10239_10383# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1556 a_9033_4399# _031_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1557 a_9390_6941# a_9117_6575# a_9305_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1558 a_4988_10933# a_4801_10973# a_4901_11191# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X1559 VPWR net10 a_9043_5487# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1560 _028_ a_8123_5487# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X1561 clknet_0_clk a_5433_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1562 VGND net12 a_9687_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1563 ones[4] a_10239_10383# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1564 VGND a_4434_9572# a_4363_9673# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X1565 VPWR a_3819_4917# net3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1566 VGND clknet_1_0__leaf_clk a_4443_4949# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1567 VPWR a_9648_2741# _045_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1568 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1569 a_5445_7439# _069_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1570 a_7350_4511# a_7182_4765# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1572 _046_ net4 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1573 a_4307_6727# a_4403_6549# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1574 a_3099_8029# a_2235_7663# a_2842_7775# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1575 VGND _073_ a_2297_7485# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1576 a_3593_8181# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1577 VGND a_5496_9269# _026_ VGND sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.143 ps=1.09 w=0.65 l=0.15
X1578 a_7987_7351# a_8083_7351# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1579 _071_ a_6835_5853# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.101875 ps=0.99 w=0.65 l=0.15
X1580 a_8231_4649# net2 _024_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1581 ones[7] a_9687_4943# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1582 a_4781_9673# a_4234_9417# a_4434_9572# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X1583 a_4807_3855# _028_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1584 VPWR a_7102_6575# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1585 a_2271_10205# a_1573_9839# a_2014_9951# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1586 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1587 _025_ a_1773_11191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1588 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1589 VGND a_4663_8029# a_4831_7931# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1590 a_9777_2767# _035_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1591 a_4035_9813# a_4326_10113# a_4277_10205# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X1592 VPWR counter\[4\] a_7843_5737# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1593 clknet_1_1__leaf_clk a_7102_6575# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1594 VGND a_5433_7637# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1595 VPWR _024_ a_2419_2767# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.26 ps=2.52 w=1 l=0.15
X1596 a_8849_10749# counter\[5\] a_8767_10749# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X1597 a_3141_4943# _011_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1598 net1 a_10199_3285# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1599 VPWR _024_ a_2734_6575# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X1600 _084_ net5 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1601 a_2253_5853# a_1915_5639# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X1602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1603 net4 a_9247_6005# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1604 VPWR a_8574_7396# a_8503_7497# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X1605 VPWR net6 a_7263_7637# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07455 ps=0.775 w=0.42 l=0.15
X1606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1607 a_6814_8207# a_6541_8213# a_6729_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1608 a_6817_6037# a_6651_6037# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1609 VPWR a_3267_7931# a_3183_8029# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1610 VPWR counter\[0\] _058_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1611 VGND clknet_1_1__leaf_clk a_8215_6037# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1612 clknet_1_1__leaf_clk a_7102_6575# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1613 a_6189_6825# _036_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1614 a_9390_8029# a_9117_7663# a_9305_7663# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1615 VGND clknet_1_1__leaf_clk a_5271_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1616 VGND a_8527_4943# a_8695_4917# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1617 a_4081_6575# counter\[4\] a_4009_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1618 a_1860_10933# a_1673_10973# a_1773_11191# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X1619 a_4319_9813# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1620 a_7607_4765# a_6743_4399# a_7350_4511# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1621 VGND a_3593_8181# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1622 a_4035_9813# a_4319_9813# a_4254_9839# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X1623 VGND a_7258_6005# a_7216_6409# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1624 VPWR a_10199_2197# net2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1625 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X1626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1627 a_4725_6397# _055_ a_4653_6397# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1628 VGND a_7833_8903# _055_ VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1629 VGND _074_ a_5731_3311# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1630 VGND a_4319_9813# a_4326_10113# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1631 a_3300_9269# _052_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1632 VPWR a_5433_7637# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1633 a_3777_5321# a_2787_4949# a_3651_4943# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1634 a_2143_7232# _072_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1635 a_4307_6727# a_4403_6549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1636 clknet_0_clk a_5433_7637# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X1637 VGND _035_ a_8013_3087# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1638 a_2431_5487# a_2295_5461# a_2011_5461# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X1639 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1640 _044_ net12 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1641 VPWR _031_ _039_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X1642 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1643 VPWR _086_ a_3851_6005# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0588 ps=0.7 w=0.42 l=0.15
X1644 VPWR a_4135_4373# _061_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27995 pd=1.615 as=0.165 ps=1.33 w=1 l=0.15
X1645 VPWR net10 _040_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1646 VGND net6 a_10239_4399# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1647 a_9122_2223# counter\[0\] a_9036_2223# VGND sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1648 VGND clknet_1_0__leaf_clk a_5547_8751# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1649 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X1650 VGND a_8971_9269# a_8929_9673# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1651 VGND a_3851_6005# _035_ VGND sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.169 ps=1.82 w=0.65 l=0.15
X1652 a_8654_6031# a_8215_6037# a_8569_6031# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1653 VPWR a_6982_8181# a_6909_8207# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1654 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1655 VPWR _051_ a_9411_7119# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1656 VPWR a_7343_7351# _063_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X1657 clknet_1_0__leaf_clk a_3593_8181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1658 a_6511_5461# counter\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X1659 VPWR a_7775_4667# a_7691_4765# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1660 VPWR _061_ a_7616_7351# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1087 ps=1.36 w=0.42 l=0.15
X1661 VGND counter\[4\] a_9963_5263# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1662 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1663 _050_ counter\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1664 a_2295_5461# clknet_1_0__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1665 a_5997_8527# counter\[7\] _073_ VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1666 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1667 _030_ a_4901_11191# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1668 _050_ a_5018_5461# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1669 a_8367_7337# clknet_1_1__leaf_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1670 VGND _035_ a_2924_6575# VGND sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X1671 a_6495_9117# a_5713_8751# a_6411_9117# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1672 a_8780_6409# a_8381_6037# a_8654_6031# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1673 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1674 VGND a_2014_9951# a_1972_9839# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1675 a_7258_6005# a_7090_6031# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1676 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1677 VGND _083_ a_4707_10703# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.095875 ps=0.945 w=0.65 l=0.15
R0 clk.n11 clk.n0 184.768
R1 clk.n10 clk.n2 184.768
R2 clk.n9 clk.n4 184.768
R3 clk.n8 clk.n6 184.768
R4 clk clk.n11 173.609
R5 clk.n11 clk.n1 146.208
R6 clk.n10 clk.n3 146.208
R7 clk.n9 clk.n5 146.208
R8 clk.n8 clk.n7 146.208
R9 clk clk.n12 56.3937
R10 clk.n11 clk.n10 40.6397
R11 clk.n10 clk.n9 40.6397
R12 clk.n9 clk.n8 40.6397
R13 clk.n12 clk 10.3624
R14 clk.n12 clk 3.45447
R15 ones[0].n0 ones[0] 79.8638
R16 ones[0] ones[0].n0 14.4176
R17 ones[0].n0 ones[0] 4.18512
R18 ones[10] ones[10].n0 83.7028
R19 ones[10].n0 ones[10] 15.9152
R20 ones[10].n0 ones[10] 0.0316459
R21 ones[1].n0 ones[1] 79.7088
R22 ones[1].n1 ones[1] 15.9152
R23 ones[1].n0 ones[1] 9.4552
R24 ones[1].n1 ones[1].n0 3.99458
R25 ones[1] ones[1].n1 0.0316459
R26 ones[2].n0 ones[2] 19.3182
R27 ones[2].n0 ones[2] 16.0107
R28 ones[2] ones[2].n0 0.030369
R29 ones[3].n0 ones[3] 79.8638
R30 ones[3].n0 ones[3] 9.4552
R31 ones[3] ones[3].n0 4.18512
R32 ones[4] ones[4].n0 1477.1
R33 ones[4].n0 ones[4] 80.894
R34 ones[4] ones[4].n1 14.114
R35 ones[4].n1 ones[4] 12.0894
R36 ones[4].n1 ones[4] 4.03013
R37 ones[4].n0 ones[4] 2.84494
R38 ones[5].n0 ones[5] 16.0107
R39 ones[5] ones[5].n0 14.2665
R40 ones[5].n0 ones[5] 0.030369
R41 ones[6].n0 ones[6] 14.5694
R42 ones[6].n0 ones[6] 12.0099
R43 ones[6] ones[6].n0 4.03013
R44 ones[7] ones[7].n0 1477.1
R45 ones[7].n0 ones[7] 80.894
R46 ones[7] ones[7].n1 14.114
R47 ones[7].n1 ones[7] 12.0894
R48 ones[7].n1 ones[7] 4.03013
R49 ones[7].n0 ones[7] 2.84494
R50 ones[8].n0 ones[8] 79.8638
R51 ones[8] ones[8].n0 18.0605
R52 ones[8].n0 ones[8] 4.18512
R53 ones[9].n0 ones[9] 18.4075
R54 ones[9].n0 ones[9] 16.0107
R55 ones[9] ones[9].n0 0.030369
R56 pulse.n2 pulse.n0 224.984
R57 pulse.n2 pulse.n1 187.714
R58 pulse pulse.n2 153.957
R59 pulse pulse.n3 10.2766
R60 pulse.n3 pulse 9.06717
R61 pulse.n3 pulse 3.02272
R62 ready.n0 ready 79.8638
R63 ready ready.n0 14.4176
R64 ready.n0 ready 4.18512
R65 rst.n2 rst.n0 224.984
R66 rst.n2 rst.n1 187.714
R67 rst.n3 rst.n2 152
R68 rst rst.n3 11.3433
R69 rst.n3 rst 1.95606
C0 counter\[1\] _028_ 0.875604f
C1 counter\[4\] _031_ 0.112206f
C2 ones[6] ones[8] 0.228608f
C3 _030_ _080_ 0.241274f
C4 _053_ _028_ 0.646754f
C5 net9 counter\[4\] 0.110581f
C6 counter\[10\] counter\[8\] 0.450807f
C7 ones[3] a_9411_8751# 0.125687f
C8 _024_ VPWR 4.28369f
C9 a_2674_9117# a_2842_8863# 0.239923f
C10 a_6099_10089# VPWR 0.185193f
C11 a_7407_8181# VPWR 0.457611f
C12 _049_ _018_ 0.260675f
C13 _021_ counter\[7\] 0.383481f
C14 a_3851_6005# VPWR 0.399487f
C15 _052_ a_3300_9269# 0.167045f
C16 counter\[6\] VPWR 2.64918f
C17 clknet_1_0__leaf_clk _017_ 0.167962f
C18 counter\[0\] _009_ 0.706492f
C19 a_8215_6037# clknet_1_1__leaf_clk 0.232623f
C20 a_8546_9269# a_7939_9301# 0.136009f
C21 _020_ a_9117_7663# 0.272277f
C22 ones[6] ones[2] 0.170254f
C23 ones[8] VPWR 0.394076f
C24 a_3651_4943# VPWR 0.194938f
C25 clk _063_ 0.111323f
C26 _086_ VPWR 3.58218f
C27 a_4687_6549# counter\[8\] 0.100618f
C28 net2 clknet_1_1__leaf_clk 0.167974f
C29 VPWR _031_ 3.1502f
C30 _080_ counter\[1\] 0.186966f
C31 ones[3] _013_ 0.275659f
C32 _053_ _060_ 0.169705f
C33 net9 VPWR 3.6191f
C34 a_5433_7637# VPWR 1.27923f
C35 clknet_0_clk counter\[8\] 0.20746f
C36 _002_ _008_ 0.639599f
C37 ones[2] VPWR 0.374056f
C38 a_1573_9839# a_2014_9951# 0.127288f
C39 _029_ _033_ 0.381626f
C40 net7 net11 0.153279f
C41 _065_ _061_ 0.280887f
C42 _015_ VPWR 0.451017f
C43 a_6817_6037# _014_ 0.174803f
C44 a_7663_4949# clknet_1_1__leaf_clk 0.226312f
C45 net3 net11 0.601931f
C46 _064_ counter\[4\] 0.370368f
C47 _048_ a_3137_4765# 0.110562f
C48 VPWR a_2511_2223# 0.220799f
C49 a_3799_8751# _026_ 0.422822f
C50 a_5437_4399# VPWR 0.300444f
C51 a_8951_7663# a_9558_7775# 0.141453f
C52 a_8083_7351# a_8374_7241# 0.189491f
C53 a_5043_4564# _015_ 0.108031f
C54 ones[2] a_10239_4399# 0.110251f
C55 clknet_1_0__leaf_clk a_3593_8181# 1.65598f
C56 a_4326_10113# VPWR 0.281484f
C57 _069_ _010_ 0.357287f
C58 _023_ _086_ 0.104651f
C59 _048_ a_8355_4074# 0.220577f
C60 a_9815_6941# a_9117_6575# 0.194916f
C61 a_7683_6005# a_7515_6031# 0.310858f
C62 _035_ clknet_1_0__leaf_clk 0.161304f
C63 a_6324_10029# VPWR 0.242368f
C64 _025_ _024_ 0.367753f
C65 _074_ VPWR 0.595788f
C66 _024_ _041_ 0.300244f
C67 _068_ VPWR 3.00196f
C68 _064_ VPWR 1.70086f
C69 a_3099_8029# VPWR 0.194219f
C70 a_6541_8213# counter\[0\] 0.114754f
C71 _070_ _053_ 0.188931f
C72 net9 a_1761_2999# 0.164804f
C73 _016_ _001_ 0.137513f
C74 _025_ _086_ 0.739186f
C75 _034_ _021_ 0.136806f
C76 a_2842_7775# VPWR 0.186717f
C77 _025_ _031_ 0.132251f
C78 a_4238_7119# VPWR 0.242589f
C79 a_6375_8213# clknet_1_1__leaf_clk 0.267046f
C80 _020_ net3 0.137057f
C81 ones[6] a_9043_5487# 0.109606f
C82 _033_ counter\[5\] 0.270548f
C83 clk rst 0.142961f
C84 _083_ net14 0.125249f
C85 _025_ net9 0.27762f
C86 _082_ VPWR 0.368581f
C87 counter\[7\] counter\[9\] 1.25284f
C88 a_6982_8181# a_6375_8213# 0.136009f
C89 ones[3] _022_ 0.151687f
C90 a_9983_6843# VPWR 0.469402f
C91 a_1915_5639# counter\[10\] 0.16559f
C92 _079_ counter\[5\] 1.33894f
C93 net5 _020_ 0.179533f
C94 a_5547_8751# a_5986_9117# 0.271965f
C95 a_1407_9839# a_1846_10205# 0.273138f
C96 counter\[7\] _076_ 0.258961f
C97 _010_ _065_ 0.432574f
C98 counter\[9\] _052_ 0.105148f
C99 a_7258_6005# VPWR 0.176757f
C100 clknet_1_0__leaf_clk net12 0.41143f
C101 counter\[0\] a_4831_7931# 0.16095f
C102 _071_ net13 0.969674f
C103 counter\[9\] _076_ 0.152223f
C104 VPWR a_8503_7497# 0.181073f
C105 clk _062_ 0.106064f
C106 a_9043_5487# VPWR 0.239898f
C107 _052_ _076_ 0.889986f
C108 ones[1] a_9503_8207# 0.123945f
C109 net4 a_7531_2741# 0.153084f
C110 a_2842_7775# a_2235_7663# 0.141453f
C111 net2 _070_ 0.194475f
C112 a_1915_5639# a_2011_5461# 0.310858f
C113 _020_ _045_ 0.11917f
C114 _027_ _010_ 0.412807f
C115 a_2502_5461# VPWR 0.25335f
C116 a_4694_6849# a_4687_6549# 0.962281f
C117 a_9735_5639# VPWR 0.199464f
C118 a_9965_11177# VPWR 0.202998f
C119 _024_ _001_ 0.166365f
C120 a_6579_9019# VPWR 0.424855f
C121 _013_ a_10103_9514# 0.108607f
C122 a_4307_6727# VPWR 0.377444f
C123 _038_ _033_ 0.598036f
C124 a_2849_5487# _010_ 0.114661f
C125 _024_ _053_ 0.612489f
C126 a_1773_11191# VPWR 0.25196f
C127 _029_ _011_ 0.212597f
C128 counter\[1\] counter\[6\] 0.501437f
C129 _038_ _079_ 0.118528f
C130 _049_ net7 0.632631f
C131 _001_ _086_ 0.193853f
C132 _083_ _028_ 0.331512f
C133 _039_ net10 0.174223f
C134 net10 _062_ 0.488358f
C135 a_8727_8181# VPWR 0.46728f
C136 _074_ a_5731_3311# 0.192864f
C137 _053_ counter\[6\] 0.392746f
C138 a_2409_4445# _024_ 0.103529f
C139 counter\[1\] _086_ 0.71637f
C140 clknet_1_0__leaf_clk _033_ 0.119941f
C141 counter\[1\] _031_ 0.352568f
C142 net6 counter\[4\] 0.357531f
C143 clknet_1_0__leaf_clk a_3799_7125# 0.226938f
C144 counter\[4\] counter\[8\] 0.680584f
C145 _053_ _031_ 0.686826f
C146 _079_ clknet_1_0__leaf_clk 0.177798f
C147 net9 counter\[1\] 0.319692f
C148 _029_ counter\[3\] 0.456819f
C149 a_6541_8213# a_7239_8207# 0.192261f
C150 _034_ counter\[7\] 0.392376f
C151 a_4981_6263# VPWR 0.142592f
C152 a_4797_4943# _006_ 0.115651f
C153 net9 _053_ 1.9697f
C154 _034_ counter\[9\] 0.793112f
C155 _020_ _054_ 1.20338f
C156 a_4609_4949# VPWR 0.284805f
C157 _069_ _049_ 0.125385f
C158 a_9558_7775# VPWR 0.184503f
C159 ones[7] net11 0.112977f
C160 net5 _009_ 0.476601f
C161 a_7843_5737# net7 0.104218f
C162 net4 VPWR 1.30325f
C163 net2 _024_ 0.3743f
C164 _063_ _061_ 0.451554f
C165 counter\[0\] clknet_1_0__leaf_clk 0.375646f
C166 _002_ net12 0.107766f
C167 _048_ VPWR 1.10875f
C168 _040_ counter\[5\] 0.418456f
C169 _053_ a_2511_2223# 0.244085f
C170 a_2401_8751# VPWR 0.306913f
C171 net6 VPWR 0.942245f
C172 _071_ net7 0.621015f
C173 a_7749_2767# VPWR 0.238674f
C174 VPWR counter\[8\] 6.17029f
C175 clknet_1_1__leaf_clk _055_ 0.365758f
C176 a_7775_4667# a_7607_4765# 0.310858f
C177 a_9983_7931# a_9815_8029# 0.310858f
C178 net8 counter\[4\] 0.34181f
C179 a_4609_4949# _006_ 0.234986f
C180 _036_ net3 0.172754f
C181 _052_ _050_ 0.182759f
C182 net2 _031_ 0.783756f
C183 _071_ net5 0.396183f
C184 a_5710_4765# VPWR 0.252597f
C185 counter\[1\] _068_ 0.132428f
C186 net6 a_10239_4399# 0.242757f
C187 net2 net9 0.102639f
C188 a_2401_7663# clknet_1_0__leaf_clk 0.474333f
C189 clk VPWR 1.10362f
C190 _064_ _053_ 0.614779f
C191 a_4526_9813# VPWR 0.240196f
C192 a_3267_7931# counter\[4\] 0.118604f
C193 _044_ counter\[8\] 0.13659f
C194 _071_ _069_ 0.226087f
C195 ones[1] _013_ 0.160999f
C196 counter\[2\] _050_ 0.214979f
C197 net10 counter\[4\] 1.02293f
C198 net9 a_10239_8751# 0.23256f
C199 net8 VPWR 3.01586f
C200 clknet_1_1__leaf_clk _051_ 0.121133f
C201 a_3847_3463# a_4120_3291# 0.167615f
C202 a_3421_3855# a_3521_3971# 0.167615f
C203 _049_ _054_ 0.22835f
C204 _067_ net11 0.12833f
C205 _086_ a_1673_10973# 0.162783f
C206 _008_ net12 0.127776f
C207 _008_ net1 0.715709f
C208 a_6060_6549# net10 0.114036f
C209 _043_ _046_ 0.125802f
C210 _080_ _055_ 0.209461f
C211 counter\[7\] net12 0.446004f
C212 counter\[7\] net1 0.281998f
C213 a_8767_10749# counter\[5\] 0.163587f
C214 _028_ _051_ 0.243308f
C215 a_3267_7931# VPWR 0.399003f
C216 a_2295_5461# clknet_1_0__leaf_clk 0.2901f
C217 _025_ net4 0.477252f
C218 a_9861_5737# a_9735_5639# 0.159564f
C219 net10 VPWR 1.80349f
C220 a_4663_7119# VPWR 0.169818f
C221 clknet_1_0__leaf_clk a_1407_9839# 0.227136f
C222 a_8075_3285# counter\[6\] 0.109662f
C223 _047_ _035_ 0.976036f
C224 _032_ VPWR 0.366191f
C225 _013_ net14 0.359497f
C226 a_3267_9019# a_3099_9117# 0.310858f
C227 _073_ _086_ 0.184068f
C228 _043_ _057_ 0.12654f
C229 net12 _003_ 0.164603f
C230 _066_ clknet_1_1__leaf_clk 0.473882f
C231 _002_ counter\[0\] 0.177634f
C232 _005_ a_6743_4399# 0.120107f
C233 _011_ clknet_1_0__leaf_clk 0.589997f
C234 a_7683_6005# VPWR 0.436775f
C235 _080_ net14 0.100857f
C236 counter\[1\] a_6579_9019# 0.132055f
C237 a_10239_10383# ones[4] 0.110247f
C238 net12 counter\[2\] 0.301446f
C239 a_8951_6575# VPWR 0.498423f
C240 net7 counter\[5\] 0.551187f
C241 _005_ counter\[4\] 0.36488f
C242 _062_ _061_ 0.100134f
C243 _073_ _015_ 0.286195f
C244 _024_ _014_ 0.156736f
C245 _010_ clknet_0_clk 0.108473f
C246 a_2674_9117# VPWR 0.24626f
C247 clknet_1_0__leaf_clk counter\[3\] 0.217299f
C248 net1 a_4225_2767# 0.135549f
C249 clknet_1_0__leaf_clk _004_ 0.178509f
C250 net5 counter\[5\] 0.27231f
C251 net8 a_8091_10615# 0.163515f
C252 clknet_0_clk net11 0.744493f
C253 _046_ VPWR 0.522708f
C254 _079_ _085_ 0.598887f
C255 net8 _025_ 0.110037f
C256 _053_ a_8727_8181# 0.105177f
C257 a_1915_5639# VPWR 0.425236f
C258 ones[0] ones[4] 0.170697f
C259 a_2734_6575# _035_ 0.129472f
C260 ones[1] _022_ 0.403959f
C261 a_4443_4949# clknet_1_0__leaf_clk 0.230418f
C262 a_4694_6849# VPWR 0.274581f
C263 _079_ counter\[7\] 0.455124f
C264 _069_ counter\[5\] 0.22447f
C265 _024_ a_2419_2767# 0.134599f
C266 _083_ counter\[6\] 0.160333f
C267 counter\[9\] a_1465_2473# 0.134849f
C268 _002_ a_6375_2767# 0.11027f
C269 _016_ _055_ 0.443319f
C270 net2 a_9735_5639# 0.152427f
C271 _037_ _055_ 0.206408f
C272 _005_ VPWR 1.63149f
C273 _032_ a_1761_2999# 0.131625f
C274 clknet_1_0__leaf_clk a_2235_8751# 0.30619f
C275 a_9687_4943# net11 0.207562f
C276 _079_ _076_ 0.185726f
C277 a_8822_6005# a_8381_6037# 0.110715f
C278 _057_ VPWR 2.37778f
C279 _039_ _000_ 0.163307f
C280 _083_ _031_ 0.11153f
C281 a_5271_8751# _033_ 0.18964f
C282 counter\[7\] counter\[0\] 0.593146f
C283 _056_ VPWR 0.349222f
C284 net4 counter\[1\] 0.183189f
C285 a_7616_7351# _061_ 0.138397f
C286 net9 _083_ 0.565725f
C287 a_5018_5461# VPWR 0.195106f
C288 _048_ counter\[1\] 0.893013f
C289 _007_ a_4326_10113# 0.181012f
C290 a_2787_4949# a_3394_4917# 0.136009f
C291 net4 _053_ 0.109205f
C292 _047_ a_2787_6031# 0.121835f
C293 counter\[1\] net6 0.171572f
C294 a_4406_8863# a_3799_8751# 0.136009f
C295 _048_ _053_ 0.132328f
C296 counter\[1\] counter\[8\] 0.218036f
C297 a_2007_7828# _042_ 0.20775f
C298 a_2014_9951# VPWR 0.232866f
C299 VPWR a_7775_4667# 0.403508f
C300 a_8017_4943# _002_ 0.114788f
C301 a_9983_7931# VPWR 0.416559f
C302 a_7833_8903# counter\[0\] 0.171631f
C303 a_9926_8181# net1 0.105103f
C304 _030_ net8 0.493067f
C305 clknet_1_0__leaf_clk a_4319_9813# 0.30159f
C306 net3 clknet_1_0__leaf_clk 0.231543f
C307 net3 a_9779_9839# 0.201899f
C308 a_5271_9295# VPWR 0.19156f
C309 _033_ _017_ 0.386093f
C310 a_3799_7663# a_3965_7663# 0.966412f
C311 _035_ net12 0.396987f
C312 _035_ net1 0.253377f
C313 a_6612_3829# VPWR 0.253171f
C314 counter\[0\] counter\[2\] 0.938797f
C315 clk counter\[1\] 0.117987f
C316 _029_ a_4589_3829# 0.12292f
C317 net5 clknet_1_0__leaf_clk 0.254914f
C318 counter\[4\] _061_ 0.979704f
C319 a_3965_7663# _000_ 0.230423f
C320 a_3965_8751# a_4663_9117# 0.192261f
C321 a_5513_10089# counter\[2\] 0.136333f
C322 _039_ net11 0.22157f
C323 a_6303_4667# net9 0.109418f
C324 _023_ _057_ 0.68311f
C325 ready net6 0.143747f
C326 ones[1] ones[8] 0.217345f
C327 a_1773_11191# a_1673_10973# 0.167615f
C328 net8 counter\[1\] 0.2245f
C329 _071_ _075_ 0.275528f
C330 net2 net6 0.113552f
C331 net8 _053_ 0.161893f
C332 counter\[5\] _078_ 1.85931f
C333 _016_ clknet_1_1__leaf_clk 0.140958f
C334 _049_ counter\[10\] 0.165434f
C335 counter\[0\] _017_ 0.816079f
C336 a_4443_4949# a_4882_4943# 0.260055f
C337 a_4609_4949# a_5050_4917# 0.127288f
C338 _085_ _040_ 2.55388f
C339 a_3799_7663# counter\[4\] 0.433307f
C340 _066_ a_7625_5461# 0.113955f
C341 _061_ VPWR 2.0538f
C342 a_8951_7663# _020_ 0.140485f
C343 counter\[7\] _040_ 1.27115f
C344 _000_ counter\[4\] 0.132055f
C345 net10 counter\[1\] 0.216317f
C346 net12 net1 0.169604f
C347 net10 _053_ 0.141143f
C348 counter\[6\] net14 0.451945f
C349 _038_ _065_ 0.341106f
C350 _034_ counter\[0\] 0.154563f
C351 _011_ _085_ 0.257668f
C352 _036_ _067_ 0.144181f
C353 a_10134_10927# _072_ 0.114695f
C354 counter\[6\] _051_ 0.167339f
C355 _019_ a_1573_9839# 0.229709f
C356 _031_ net14 0.52284f
C357 a_6411_9117# a_6579_9019# 0.310858f
C358 _039_ _020_ 0.12729f
C359 _013_ _022_ 0.163537f
C360 _013_ a_8374_7241# 0.184263f
C361 _086_ _051_ 0.32257f
C362 a_3799_7663# VPWR 0.438944f
C363 net2 net8 0.142942f
C364 a_6729_8207# _008_ 0.114852f
C365 _009_ _042_ 0.13669f
C366 net7 _026_ 0.199788f
C367 _031_ _051_ 0.254741f
C368 _038_ _027_ 0.182173f
C369 _000_ VPWR 0.430233f
C370 a_9687_8751# net12 0.257694f
C371 net9 _051_ 0.101631f
C372 clknet_0_clk _009_ 0.154576f
C373 counter\[0\] _050_ 0.319973f
C374 counter\[2\] net13 0.11425f
C375 _010_ counter\[4\] 0.293578f
C376 counter\[7\] _004_ 0.205148f
C377 _024_ clknet_1_1__leaf_clk 0.746479f
C378 a_3137_4765# _049_ 0.173338f
C379 clknet_1_0__leaf_clk _054_ 0.422119f
C380 _074_ _055_ 0.185026f
C381 counter\[4\] net11 0.188475f
C382 _027_ clknet_1_0__leaf_clk 0.109659f
C383 a_3521_3971# VPWR 0.205438f
C384 _018_ _050_ 0.663593f
C385 clknet_1_1__leaf_clk counter\[6\] 0.111415f
C386 clknet_1_0__leaf_clk _078_ 0.147325f
C387 _073_ counter\[8\] 0.333428f
C388 a_5625_4399# _016_ 0.120612f
C389 a_9117_6575# _018_ 0.278513f
C390 clknet_1_1__leaf_clk _086_ 0.385842f
C391 _047_ _040_ 0.173723f
C392 _069_ _002_ 0.767788f
C393 _003_ _004_ 0.486077f
C394 a_3099_9117# VPWR 0.191336f
C395 a_7090_6031# a_6651_6037# 0.259867f
C396 a_7258_6005# a_6817_6037# 0.110715f
C397 ones[4] _031_ 0.143222f
C398 counter\[6\] _028_ 0.480888f
C399 _079_ net1 1.22417f
C400 a_6909_4399# a_7607_4765# 0.192341f
C401 counter\[3\] counter\[2\] 0.512581f
C402 _010_ VPWR 2.24831f
C403 _059_ a_2511_2223# 0.204282f
C404 _043_ _020_ 0.909789f
C405 VPWR net11 3.58797f
C406 a_4238_8029# a_3799_7663# 0.260055f
C407 a_4406_7775# a_3965_7663# 0.117154f
C408 _081_ _016_ 0.21448f
C409 counter\[0\] a_5713_8751# 0.455193f
C410 _005_ a_5823_7119# 0.107307f
C411 _057_ _053_ 0.202778f
C412 _068_ _051_ 0.157282f
C413 _015_ clknet_1_1__leaf_clk 0.134723f
C414 a_4443_4949# counter\[2\] 0.311046f
C415 ones[5] VPWR 0.516632f
C416 net4 _014_ 0.112062f
C417 _008_ net7 0.159054f
C418 _039_ _049_ 0.23294f
C419 a_5437_4399# clknet_1_1__leaf_clk 0.452985f
C420 _003_ a_2235_8751# 0.250656f
C421 a_1573_9839# a_2271_10205# 0.196846f
C422 counter\[0\] net12 0.941195f
C423 net3 _085_ 0.198804f
C424 counter\[3\] _017_ 0.191384f
C425 net4 _083_ 0.101239f
C426 _014_ counter\[8\] 0.34718f
C427 a_2051_4943# VPWR 0.286902f
C428 _020_ counter\[4\] 0.107719f
C429 net5 _085_ 0.100679f
C430 _049_ a_3203_7351# 0.135886f
C431 _040_ _050_ 0.102709f
C432 net3 _052_ 0.888921f
C433 net7 _076_ 0.231435f
C434 a_8367_7337# a_8574_7396# 0.260055f
C435 a_4135_4373# VPWR 0.497606f
C436 net3 _076_ 0.222839f
C437 _074_ clknet_1_1__leaf_clk 0.220726f
C438 a_10136_4943# VPWR 0.257702f
C439 VPWR a_9963_4399# 0.269603f
C440 _035_ net13 0.111845f
C441 net5 _052_ 0.804571f
C442 _069_ counter\[7\] 1.44016f
C443 _034_ _004_ 1.18836f
C444 net5 _076_ 0.307118f
C445 net7 counter\[2\] 0.701177f
C446 _011_ _050_ 0.132742f
C447 _069_ counter\[9\] 0.992988f
C448 a_2007_7828# VPWR 0.255977f
C449 net3 counter\[2\] 1.46437f
C450 clk _083_ 0.160568f
C451 a_8822_6005# VPWR 0.181132f
C452 _020_ VPWR 1.40428f
C453 a_9735_5639# net14 0.14297f
C454 net8 _014_ 0.309619f
C455 _072_ _019_ 0.838435f
C456 a_2776_7119# VPWR 0.235994f
C457 counter\[0\] _033_ 0.113183f
C458 _011_ a_2953_4949# 0.562122f
C459 counter\[1\] _061_ 0.807381f
C460 _077_ _075_ 0.257784f
C461 a_4406_7775# VPWR 0.180791f
C462 net8 _083_ 3.59944f
C463 counter\[3\] _050_ 0.484857f
C464 net4 a_6817_6037# 0.457319f
C465 a_4227_9513# VPWR 0.640169f
C466 net5 a_4831_9019# 0.105942f
C467 _053_ _061_ 0.495569f
C468 net7 _017_ 0.11f
C469 _069_ counter\[2\] 0.280393f
C470 net12 _040_ 0.171764f
C471 _029_ _039_ 0.100116f
C472 net1 _040_ 0.20993f
C473 _024_ _016_ 0.137566f
C474 _049_ counter\[4\] 0.27884f
C475 a_8822_6005# a_8654_6031# 0.239923f
C476 net12 net13 0.520804f
C477 net1 net13 0.565713f
C478 a_5871_9527# VPWR 0.210399f
C479 net10 _083_ 0.205287f
C480 a_6743_4399# a_6909_4399# 0.959715f
C481 _037_ counter\[6\] 0.484043f
C482 _012_ clknet_1_0__leaf_clk 0.6349f
C483 counter\[9\] _065_ 0.109199f
C484 a_4406_7093# a_3799_7125# 0.136009f
C485 a_3965_7125# _015_ 0.561623f
C486 _022_ _086_ 2.09057f
C487 _009_ counter\[4\] 0.856303f
C488 counter\[7\] _054_ 0.672638f
C489 _069_ _047_ 0.347614f
C490 a_2787_6031# _040_ 0.116577f
C491 clknet_1_0__leaf_clk _063_ 0.150636f
C492 net9 _022_ 0.67748f
C493 _027_ counter\[7\] 0.122005f
C494 _082_ _080_ 1.09563f
C495 _085_ _078_ 0.407763f
C496 _049_ VPWR 1.0681f
C497 _052_ _054_ 0.337117f
C498 _027_ counter\[9\] 0.351694f
C499 counter\[7\] _078_ 0.973563f
C500 a_4406_7775# a_4238_8029# 0.239923f
C501 VPWR a_8268_2741# 0.180986f
C502 a_4227_9513# a_4234_9417# 0.970213f
C503 a_7987_7351# VPWR 0.395272f
C504 _053_ a_3521_3971# 0.100942f
C505 _081_ _074_ 0.202171f
C506 net3 _050_ 0.373241f
C507 _048_ _051_ 0.189355f
C508 net6 _051_ 0.35513f
C509 a_5437_4399# _016_ 0.194614f
C510 _035_ net3 0.202475f
C511 a_4901_11191# VPWR 0.206793f
C512 _071_ counter\[4\] 0.142807f
C513 a_4801_10973# a_4901_11191# 0.167615f
C514 _076_ _078_ 0.302306f
C515 _009_ VPWR 2.1475f
C516 a_10134_10927# VPWR 0.217556f
C517 clknet_1_0__leaf_clk _042_ 0.325897f
C518 a_6979_10901# _071_ 0.168913f
C519 _010_ counter\[1\] 0.262662f
C520 a_7939_9301# net7 0.423465f
C521 a_7102_6575# net11 0.220052f
C522 VPWR a_6909_4399# 0.320082f
C523 ones[6] _071_ 0.100567f
C524 _049_ _006_ 0.614372f
C525 counter\[1\] net11 1.00294f
C526 _014_ _005_ 0.547735f
C527 a_7263_7637# net1 0.132942f
C528 a_7843_5737# VPWR 0.210702f
C529 _053_ net11 0.226832f
C530 _024_ _086_ 1.58345f
C531 _016_ _074_ 0.225695f
C532 net4 clknet_1_1__leaf_clk 0.591612f
C533 a_5547_8751# VPWR 0.598327f
C534 _069_ _035_ 0.230519f
C535 a_6060_6549# _036_ 0.148634f
C536 _024_ _031_ 0.763267f
C537 VPWR a_1846_10205# 0.293883f
C538 _011_ _079_ 0.832112f
C539 net6 clknet_1_1__leaf_clk 0.485145f
C540 a_5871_9527# _041_ 0.201967f
C541 _071_ VPWR 2.6663f
C542 ones[3] ones[5] 0.123415f
C543 _035_ _045_ 0.842383f
C544 _024_ net9 0.584321f
C545 _021_ a_8381_6037# 0.255478f
C546 clknet_1_1__leaf_clk counter\[8\] 0.112433f
C547 counter\[6\] _031_ 0.498101f
C548 net8 _051_ 0.218484f
C549 _036_ VPWR 0.28636f
C550 net4 _028_ 0.624754f
C551 net9 counter\[6\] 0.317728f
C552 net7 net12 0.41731f
C553 _086_ _031_ 0.248361f
C554 a_3847_6727# VPWR 0.182946f
C555 a_4135_4373# counter\[1\] 0.169857f
C556 net3 net12 0.139261f
C557 net3 net1 0.735136f
C558 _011_ counter\[0\] 0.191378f
C559 _082_ _016_ 0.511494f
C560 net9 _086_ 0.236918f
C561 _009_ a_4234_9417# 0.261284f
C562 net9 _031_ 0.265824f
C563 a_10136_4943# _053_ 0.209447f
C564 clk clknet_1_1__leaf_clk 0.149771f
C565 net10 net14 0.185922f
C566 _029_ VPWR 0.896414f
C567 net5 net12 0.681877f
C568 net5 net1 0.763374f
C569 a_8105_9301# VPWR 0.293336f
C570 _038_ _039_ 0.124421f
C571 ones[2] _031_ 0.362981f
C572 _034_ _027_ 1.65938f
C573 a_8374_7241# a_8503_7497# 0.11316f
C574 _065_ _050_ 0.229426f
C575 a_6541_8213# VPWR 0.309888f
C576 counter\[0\] counter\[3\] 0.24495f
C577 net8 clknet_1_1__leaf_clk 0.310308f
C578 _058_ counter\[7\] 0.146423f
C579 _020_ _053_ 0.448211f
C580 _035_ _065_ 0.821095f
C581 _024_ _074_ 0.414883f
C582 counter\[3\] a_5513_10089# 0.126519f
C583 net8 a_10239_10383# 0.233688f
C584 _039_ clknet_1_0__leaf_clk 0.373831f
C585 a_3819_4917# net3 0.145863f
C586 a_8527_4943# a_7829_4949# 0.192261f
C587 a_3476_7351# counter\[8\] 0.116646f
C588 net12 _045_ 0.710507f
C589 net1 _045_ 0.746281f
C590 ones[5] a_10239_8751# 0.110675f
C591 a_8102_4943# VPWR 0.241556f
C592 ready a_9963_4399# 0.110391f
C593 _068_ counter\[6\] 0.137306f
C594 _075_ _076_ 0.173078f
C595 _027_ _050_ 0.131492f
C596 counter\[5\] counter\[4\] 0.973378f
C597 _064_ counter\[6\] 0.220033f
C598 a_10199_3285# net1 0.173518f
C599 _005_ _055_ 0.109819f
C600 a_9247_6005# VPWR 0.388515f
C601 _002_ a_7829_4949# 0.253372f
C602 counter\[7\] _067_ 0.221012f
C603 a_7987_7351# a_8083_7351# 0.310858f
C604 net10 clknet_1_1__leaf_clk 0.318041f
C605 net3 _033_ 0.102226f
C606 a_5271_4399# a_5878_4511# 0.136009f
C607 a_2401_7663# _004_ 0.213056f
C608 _056_ _055_ 0.109815f
C609 _071_ _025_ 1.25264f
C610 _012_ _085_ 0.126073f
C611 _082_ _024_ 0.207777f
C612 _058_ counter\[2\] 0.469074f
C613 a_4831_7931# VPWR 0.426797f
C614 a_4434_9572# VPWR 0.251798f
C615 a_8822_6005# a_8215_6037# 0.136009f
C616 a_7711_3463# counter\[4\] 0.196841f
C617 a_7683_6005# clknet_1_1__leaf_clk 0.10999f
C618 _030_ a_4901_11191# 0.103764f
C619 a_8270_4917# a_8102_4943# 0.239923f
C620 counter\[7\] _063_ 0.11002f
C621 _010_ _073_ 0.921717f
C622 counter\[5\] VPWR 2.66496f
C623 a_8951_6575# clknet_1_1__leaf_clk 0.22115f
C624 counter\[7\] counter\[10\] 0.274231f
C625 a_8546_9269# VPWR 0.189552f
C626 counter\[9\] counter\[10\] 0.919353f
C627 _010_ a_6375_8213# 0.463367f
C628 _019_ VPWR 0.804658f
C629 counter\[0\] net3 0.482611f
C630 _037_ a_4981_6263# 0.105515f
C631 _072_ counter\[7\] 1.39989f
C632 _043_ clknet_1_0__leaf_clk 0.44364f
C633 a_6909_4399# a_7350_4511# 0.112272f
C634 a_6743_4399# a_7182_4765# 0.260055f
C635 _012_ _003_ 0.184188f
C636 net1 _054_ 0.667402f
C637 _069_ a_1465_2473# 0.123428f
C638 net7 _018_ 0.634217f
C639 net5 counter\[0\] 0.213603f
C640 a_7711_3463# VPWR 0.345046f
C641 _044_ counter\[5\] 0.157403f
C642 a_4694_6849# clknet_1_1__leaf_clk 0.376909f
C643 a_7616_7351# a_7343_7351# 0.167615f
C644 _064_ a_6324_10029# 0.201417f
C645 _068_ _064_ 0.982966f
C646 a_9122_2223# VPWR 0.199942f
C647 _069_ counter\[0\] 0.418151f
C648 clknet_1_0__leaf_clk counter\[4\] 0.168726f
C649 _039_ _026_ 0.869945f
C650 _024_ a_1773_11191# 0.20318f
C651 _052_ _042_ 0.595131f
C652 a_4227_9513# a_4363_9673# 0.141453f
C653 _005_ clknet_1_1__leaf_clk 0.38254f
C654 _014_ _010_ 0.13484f
C655 a_9551_9527# VPWR 0.197306f
C656 _066_ _005_ 0.448496f
C657 a_2409_5263# counter\[9\] 0.101438f
C658 _061_ _055_ 0.43733f
C659 a_5496_9269# _026_ 0.145227f
C660 _038_ VPWR 1.34534f
C661 _056_ clknet_1_1__leaf_clk 0.956141f
C662 _003_ _042_ 0.198494f
C663 _033_ _065_ 0.204933f
C664 _030_ _029_ 1.11415f
C665 a_10199_3285# pulse 0.226298f
C666 VPWR a_7182_4765# 0.265764f
C667 _083_ net11 0.102894f
C668 net2 _049_ 0.196598f
C669 a_9687_10927# net13 0.215507f
C670 a_8123_5487# net7 0.157979f
C671 a_9815_6941# VPWR 0.187585f
C672 a_8123_5487# net3 0.114389f
C673 clknet_1_0__leaf_clk VPWR 4.19422f
C674 a_9779_9839# VPWR 0.232349f
C675 _077_ VPWR 1.15656f
C676 net8 _016_ 0.466971f
C677 ones[7] net1 0.155178f
C678 net7 _040_ 0.246539f
C679 a_3965_7125# a_4663_7119# 0.191992f
C680 VPWR a_2271_10205# 0.204828f
C681 _000_ a_2879_8207# 0.109088f
C682 a_3943_9527# VPWR 0.185352f
C683 _029_ counter\[1\] 0.528435f
C684 net3 net13 1.30775f
C685 _079_ _078_ 0.164385f
C686 a_9117_7663# net3 0.166731f
C687 clknet_0_clk _017_ 0.671382f
C688 ones[9] a_9687_10927# 0.10957f
C689 a_7343_7351# VPWR 0.208185f
C690 clknet_1_0__leaf_clk _006_ 0.512896f
C691 _044_ clknet_1_0__leaf_clk 0.215043f
C692 a_6335_5461# VPWR 0.168818f
C693 a_7407_8181# counter\[8\] 0.125622f
C694 net5 net13 0.13993f
C695 clknet_1_0__leaf_clk a_2235_7663# 0.313183f
C696 counter\[6\] counter\[8\] 0.896443f
C697 a_2509_4663# VPWR 0.211641f
C698 net6 _086_ 0.166746f
C699 net4 net9 0.203703f
C700 net6 _031_ 0.158942f
C701 _039_ counter\[9\] 0.211847f
C702 _086_ counter\[8\] 0.47191f
C703 a_4687_6549# a_4823_6575# 0.136001f
C704 _048_ net9 0.599992f
C705 _023_ clknet_1_0__leaf_clk 0.113511f
C706 a_9558_6687# a_8951_6575# 0.14092f
C707 counter\[8\] _031_ 0.757795f
C708 a_3300_9269# VPWR 0.264055f
C709 _014_ a_2776_7119# 0.104948f
C710 _035_ counter\[10\] 0.224916f
C711 counter\[4\] _026_ 0.152017f
C712 clknet_1_1__leaf_clk _061_ 0.819368f
C713 net3 counter\[3\] 0.313119f
C714 _020_ a_9305_7663# 0.115579f
C715 net9 counter\[8\] 0.277893f
C716 _002_ counter\[4\] 0.107365f
C717 clk counter\[6\] 0.185443f
C718 _021_ VPWR 0.511033f
C719 counter\[9\] a_3203_7351# 0.225962f
C720 _039_ _003_ 0.102598f
C721 _055_ net11 0.36656f
C722 a_6651_6037# VPWR 0.474411f
C723 _015_ counter\[8\] 0.339981f
C724 a_2589_7663# _004_ 0.118037f
C725 _067_ net1 0.987729f
C726 a_3943_9527# a_4234_9417# 0.194892f
C727 net8 counter\[6\] 0.96701f
C728 a_8527_4943# VPWR 0.18128f
C729 clknet_0_clk a_3593_8181# 0.316596f
C730 clk a_5433_7637# 0.315386f
C731 _069_ ones[9] 0.187618f
C732 net8 _086_ 0.181359f
C733 a_2295_5461# a_2431_5487# 0.141453f
C734 _026_ VPWR 1.69281f
C735 counter\[1\] counter\[5\] 0.365458f
C736 _084_ _019_ 0.195774f
C737 _019_ _001_ 0.273075f
C738 net8 _031_ 4.8238f
C739 _070_ _057_ 0.134894f
C740 _002_ VPWR 0.563296f
C741 a_4882_4943# VPWR 0.240131f
C742 _048_ _068_ 0.122759f
C743 net8 net9 1.47097f
C744 net14 net11 0.200731f
C745 net5 a_7263_7637# 0.22043f
C746 _039_ _017_ 0.103823f
C747 _063_ net12 0.152816f
C748 a_3851_6005# net10 0.164667f
C749 net10 counter\[6\] 0.379499f
C750 _051_ net11 0.64785f
C751 a_5503_11092# _038_ 0.200768f
C752 net8 _015_ 0.395843f
C753 _014_ _049_ 0.286087f
C754 a_4601_5737# a_4351_5737# 0.144824f
C755 _008_ counter\[4\] 0.386913f
C756 net3 net7 0.360564f
C757 a_8971_9269# VPWR 0.407726f
C758 _085_ counter\[4\] 0.225183f
C759 net10 _031_ 0.216951f
C760 _079_ _075_ 0.104946f
C761 _066_ a_3521_3971# 0.200974f
C762 a_9247_6005# a_9079_6031# 0.310858f
C763 counter\[7\] counter\[4\] 0.536222f
C764 _083_ a_8268_2741# 0.133959f
C765 a_7350_4511# a_7182_4765# 0.239923f
C766 a_8102_4943# a_7663_4949# 0.260055f
C767 net5 net7 0.271187f
C768 _032_ net9 0.14175f
C769 net5 net3 2.27782f
C770 a_8951_6575# _086_ 0.356695f
C771 net2 counter\[5\] 0.146736f
C772 clknet_1_1__leaf_clk net11 1.4471f
C773 a_9011_3285# VPWR 0.461817f
C774 a_9963_4399# net14 0.220715f
C775 _058_ counter\[0\] 0.149192f
C776 _069_ net7 0.261218f
C777 net8 _074_ 0.347358f
C778 _069_ net3 0.371215f
C779 a_2971_4399# _049_ 0.12513f
C780 a_1559_2473# VPWR 0.207919f
C781 _008_ VPWR 0.982338f
C782 _047_ a_7531_2741# 0.140635f
C783 a_2589_8751# _003_ 0.123343f
C784 _085_ VPWR 1.13654f
C785 _084_ clknet_1_0__leaf_clk 0.475906f
C786 clknet_1_0__leaf_clk _001_ 0.34908f
C787 a_4831_7931# a_4663_8029# 0.310858f
C788 a_1573_9839# a_1407_9839# 0.974409f
C789 net3 _045_ 0.234448f
C790 counter\[7\] VPWR 3.36658f
C791 _058_ _018_ 0.108294f
C792 a_4434_9572# a_4363_9673# 0.239923f
C793 counter\[4\] counter\[2\] 0.269736f
C794 _027_ counter\[3\] 1.55545f
C795 _039_ _035_ 0.343623f
C796 _024_ _005_ 0.21886f
C797 a_7005_6031# _014_ 0.133039f
C798 counter\[9\] VPWR 1.3638f
C799 _047_ _043_ 1.10839f
C800 _024_ _057_ 0.108209f
C801 a_6541_8213# a_6375_8213# 0.96217f
C802 a_7108_5737# VPWR 0.195311f
C803 clknet_1_0__leaf_clk _053_ 0.126662f
C804 a_2439_10107# a_2271_10205# 0.310858f
C805 a_3267_7931# a_3099_8029# 0.310858f
C806 _052_ VPWR 0.570079f
C807 _036_ _014_ 0.116159f
C808 a_4609_4949# a_4797_4943# 0.101638f
C809 net10 _068_ 0.116128f
C810 a_3799_8751# VPWR 0.438415f
C811 net10 _064_ 0.110243f
C812 _076_ VPWR 0.893794f
C813 a_7833_8903# VPWR 0.174915f
C814 _057_ counter\[6\] 0.195928f
C815 ones[7] net13 0.136832f
C816 VPWR a_9739_6005# 0.405629f
C817 a_3847_9527# a_3943_9527# 0.310858f
C818 _003_ VPWR 1.18877f
C819 ones[0] ones[5] 0.127204f
C820 ones[1] _049_ 0.300154f
C821 _037_ _061_ 0.660469f
C822 a_5271_8751# VPWR 0.191682f
C823 a_8546_9269# a_8378_9295# 0.239923f
C824 counter\[2\] VPWR 4.3923f
C825 counter\[0\] _063_ 0.434052f
C826 _021_ a_8569_6031# 0.11532f
C827 net2 _038_ 0.129496f
C828 a_6335_5461# _053_ 0.271441f
C829 a_4831_9019# VPWR 0.372461f
C830 a_9411_7119# _049_ 0.131453f
C831 VPWR a_4225_2767# 0.242287f
C832 _073_ counter\[5\] 0.21653f
C833 net7 _054_ 0.257218f
C834 _034_ counter\[4\] 0.86423f
C835 VPWR a_8397_2767# 0.191962f
C836 a_2409_5263# _079_ 0.139107f
C837 a_3300_9269# _053_ 0.156786f
C838 _027_ net7 0.224358f
C839 a_2409_4445# a_2509_4663# 0.167615f
C840 _017_ VPWR 0.54274f
C841 a_4120_3291# VPWR 0.160005f
C842 a_9043_5487# net10 0.189002f
C843 _075_ net13 0.115905f
C844 _047_ VPWR 1.12743f
C845 _052_ a_4234_9417# 0.259739f
C846 _069_ _065_ 0.137229f
C847 _025_ counter\[7\] 0.381649f
C848 counter\[7\] _041_ 0.588032f
C849 a_2235_8751# a_2842_8863# 0.141453f
C850 a_6135_4765# VPWR 0.169772f
C851 a_7711_3463# a_8075_3285# 0.124682f
C852 _034_ VPWR 1.18289f
C853 a_5731_3311# _008_ 0.108513f
C854 a_4823_6575# VPWR 0.174392f
C855 a_3847_3463# VPWR 0.206327f
C856 counter\[6\] _061_ 0.36976f
C857 clk net4 1.38189f
C858 _002_ _053_ 0.560283f
C859 _061_ _086_ 0.371139f
C860 a_8215_6037# _021_ 0.114598f
C861 a_9926_8181# VPWR 0.189938f
C862 _083_ counter\[5\] 0.608407f
C863 a_3593_8181# VPWR 1.23f
C864 _022_ net11 0.646678f
C865 _047_ _023_ 0.175983f
C866 VPWR _050_ 1.43382f
C867 a_2734_6575# VPWR 0.445476f
C868 net8 net4 0.255551f
C869 _035_ VPWR 2.1093f
C870 a_5307_4943# VPWR 0.171286f
C871 _030_ _085_ 0.128164f
C872 a_2302_5761# _010_ 0.227178f
C873 net8 _048_ 0.111328f
C874 a_9117_6575# VPWR 0.305507f
C875 _068_ a_6612_3829# 0.185734f
C876 clknet_1_0__leaf_clk _073_ 0.111907f
C877 a_4981_6263# net10 0.193932f
C878 pulse rst 0.135916f
C879 a_7939_9301# VPWR 0.45178f
C880 a_2953_4949# VPWR 0.283391f
C881 VPWR a_8367_7337# 0.413943f
C882 clknet_1_1__leaf_clk a_6909_4399# 0.367861f
C883 a_6835_5853# VPWR 0.232606f
C884 _025_ _017_ 0.143109f
C885 net12 counter\[4\] 1.30459f
C886 a_8695_4917# a_8527_4943# 0.310858f
C887 net1 counter\[4\] 0.793814f
C888 _012_ counter\[3\] 0.278601f
C889 _043_ a_2787_6031# 0.100657f
C890 _084_ _085_ 0.125941f
C891 _085_ _001_ 0.775646f
C892 a_4319_9813# a_4455_9839# 0.136009f
C893 _027_ _065_ 0.321832f
C894 _035_ _006_ 0.573729f
C895 _007_ a_4873_9839# 0.114653f
C896 counter\[7\] _001_ 0.199605f
C897 a_8803_9295# a_8105_9301# 0.192261f
C898 _007_ clknet_1_0__leaf_clk 0.183945f
C899 _070_ _020_ 0.302608f
C900 a_6060_6549# net12 0.1351f
C901 counter\[7\] counter\[1\] 0.487933f
C902 _008_ _053_ 0.335004f
C903 _034_ a_8091_10615# 0.112526f
C904 net10 counter\[8\] 0.536843f
C905 a_5713_8751# VPWR 0.276778f
C906 _085_ _053_ 0.12899f
C907 a_4351_5737# counter\[3\] 0.141854f
C908 net3 _075_ 0.257647f
C909 _074_ _061_ 1.01237f
C910 counter\[7\] _053_ 0.314743f
C911 _068_ _061_ 0.140407f
C912 _054_ _078_ 0.135712f
C913 _064_ _061_ 0.152926f
C914 _023_ _035_ 0.279192f
C915 a_7663_4949# _002_ 0.110977f
C916 counter\[9\] _053_ 0.217527f
C917 a_5050_4917# a_4882_4943# 0.239923f
C918 _014_ clknet_1_0__leaf_clk 0.337215f
C919 _027_ _078_ 0.142745f
C920 a_4601_5737# VPWR 0.184621f
C921 net12 VPWR 2.45198f
C922 net1 VPWR 2.18353f
C923 _037_ _020_ 0.114197f
C924 a_7833_8903# counter\[1\] 0.118091f
C925 counter\[3\] _042_ 0.699761f
C926 _004_ _042_ 0.934811f
C927 a_5503_11092# _017_ 0.112747f
C928 _010_ _086_ 0.140293f
C929 a_2971_4399# _038_ 0.119667f
C930 _030_ _017_ 0.264341f
C931 _029_ clknet_1_1__leaf_clk 0.371307f
C932 _036_ _028_ 0.570599f
C933 _086_ net11 0.791436f
C934 counter\[1\] counter\[2\] 0.62994f
C935 a_9117_7663# a_9815_8029# 0.194972f
C936 _031_ net11 0.145476f
C937 net8 net10 0.339199f
C938 _053_ counter\[2\] 0.432856f
C939 a_6814_8207# VPWR 0.260461f
C940 _044_ net12 0.257227f
C941 a_2787_6031# VPWR 0.616523f
C942 a_9687_8751# VPWR 0.201839f
C943 a_6541_8213# clknet_1_1__leaf_clk 0.188445f
C944 a_8951_7663# a_9117_7663# 0.970312f
C945 a_3819_4917# VPWR 0.46711f
C946 net2 counter\[7\] 0.122145f
C947 ones[5] net9 0.204931f
C948 _073_ _026_ 0.156739f
C949 a_8231_4649# VPWR 0.350546f
C950 _063_ a_4319_9813# 0.421054f
C951 _069_ _067_ 0.53155f
C952 a_6541_8213# a_6982_8181# 0.118966f
C953 _039_ _040_ 0.217312f
C954 net2 _052_ 0.188887f
C955 _070_ _049_ 0.254557f
C956 _033_ VPWR 0.796808f
C957 counter\[0\] counter\[4\] 0.126842f
C958 a_1775_4399# VPWR 0.254009f
C959 _035_ a_9648_2741# 0.131994f
C960 a_4319_2767# VPWR 0.20096f
C961 a_6335_5461# a_6511_5461# 0.185422f
C962 a_3799_7125# VPWR 0.411253f
C963 _056_ counter\[8\] 0.696159f
C964 _079_ VPWR 0.695815f
C965 net7 _042_ 0.128769f
C966 VPWR a_1465_2473# 0.239992f
C967 _020_ counter\[6\] 0.136931f
C968 a_5271_4399# VPWR 0.41634f
C969 net2 counter\[2\] 0.498651f
C970 _037_ _049_ 0.206097f
C971 _034_ counter\[1\] 0.747626f
C972 _074_ net11 0.51498f
C973 a_7711_3463# _051_ 0.111517f
C974 a_8695_4917# counter\[2\] 0.129366f
C975 net3 clknet_0_clk 0.370845f
C976 _069_ _072_ 2.04001f
C977 a_4406_8863# VPWR 0.177439f
C978 clknet_1_1__leaf_clk counter\[5\] 0.279813f
C979 a_4153_7663# a_3965_7663# 0.101638f
C980 net2 a_4225_2767# 0.130972f
C981 counter\[0\] VPWR 2.29289f
C982 net5 clknet_0_clk 0.216045f
C983 _062_ _004_ 0.108622f
C984 _027_ _075_ 0.239202f
C985 a_7663_4949# counter\[2\] 0.424234f
C986 _058_ _027_ 0.103203f
C987 VPWR pulse 0.137491f
C988 a_5513_10089# VPWR 0.143288f
C989 a_4035_9813# VPWR 0.167017f
C990 _024_ a_5871_9527# 0.253426f
C991 _046_ net10 0.521903f
C992 counter\[1\] _050_ 0.141291f
C993 _038_ _051_ 0.10598f
C994 _043_ _040_ 0.187037f
C995 _018_ VPWR 1.08549f
C996 a_2787_4949# clknet_1_0__leaf_clk 0.314082f
C997 a_7987_7828# _009_ 0.108485f
C998 counter\[7\] _073_ 0.122441f
C999 counter\[7\] a_8075_3285# 0.280169f
C1000 _053_ _050_ 0.258014f
C1001 a_9122_2223# _059_ 0.170218f
C1002 a_6375_8213# _008_ 0.130626f
C1003 _043_ net13 0.242386f
C1004 counter\[9\] _073_ 1.05985f
C1005 a_9983_6843# net11 0.15198f
C1006 _071_ _022_ 1.51183f
C1007 a_3421_3855# _065_ 0.154412f
C1008 a_10136_4943# _064_ 0.150447f
C1009 a_2401_7663# VPWR 0.310323f
C1010 _073_ _052_ 0.124147f
C1011 a_4406_7093# VPWR 0.174364f
C1012 net4 _061_ 0.13983f
C1013 _057_ net10 0.141729f
C1014 a_2409_4445# _035_ 0.124357f
C1015 _048_ _061_ 0.18673f
C1016 a_6651_6037# a_6817_6037# 0.961627f
C1017 net6 _061_ 0.818543f
C1018 _040_ counter\[4\] 0.118924f
C1019 _056_ net10 0.111556f
C1020 a_6835_5853# _053_ 0.228449f
C1021 _007_ counter\[7\] 0.739582f
C1022 a_9390_6941# VPWR 0.243854f
C1023 _061_ counter\[8\] 0.534818f
C1024 _001_ a_5713_8751# 0.186639f
C1025 net5 a_8951_7663# 0.154621f
C1026 a_5547_8751# a_6154_8863# 0.136001f
C1027 VPWR a_6375_2767# 0.276508f
C1028 a_4901_11191# _024_ 0.243407f
C1029 a_3226_4943# VPWR 0.256946f
C1030 _027_ counter\[10\] 0.118887f
C1031 VPWR a_8574_7396# 0.257963f
C1032 a_8123_5487# VPWR 0.389503f
C1033 _022_ a_8105_9301# 0.564016f
C1034 _014_ counter\[7\] 0.367916f
C1035 counter\[10\] _078_ 0.102091f
C1036 a_2401_7663# a_2235_7663# 0.966391f
C1037 net12 a_2439_10107# 0.129063f
C1038 clk _061_ 0.460807f
C1039 counter\[1\] net12 0.177394f
C1040 a_2295_5461# VPWR 0.696157f
C1041 _077_ clknet_1_1__leaf_clk 0.422615f
C1042 _040_ VPWR 2.16885f
C1043 counter\[7\] _083_ 0.413894f
C1044 net12 _053_ 0.601855f
C1045 net1 _053_ 0.22611f
C1046 a_1407_9839# VPWR 0.756948f
C1047 _007_ counter\[2\] 0.108446f
C1048 _014_ _076_ 0.155378f
C1049 a_5986_9117# VPWR 0.255161f
C1050 a_10103_9991# _076_ 0.202345f
C1051 VPWR net13 2.01646f
C1052 _046_ _057_ 0.369408f
C1053 _004_ counter\[4\] 0.226011f
C1054 net8 _061_ 0.442481f
C1055 a_9117_7663# VPWR 0.311819f
C1056 _069_ _039_ 0.172473f
C1057 ones[9] ones[10] 0.199863f
C1058 a_3799_8751# a_4238_9117# 0.260055f
C1059 _011_ VPWR 0.265899f
C1060 _024_ _036_ 0.348547f
C1061 _039_ _045_ 0.206085f
C1062 _003_ a_3479_10004# 0.107854f
C1063 _071_ ones[8] 0.824493f
C1064 a_7239_8207# VPWR 0.191342f
C1065 _058_ _075_ 1.42232f
C1066 a_8767_10749# counter\[4\] 0.173697f
C1067 ready net1 0.20058f
C1068 ones[0] a_9779_9839# 0.110372f
C1069 ones[0] _077_ 0.207691f
C1070 _044_ net13 0.129516f
C1071 _071_ _031_ 0.391362f
C1072 ones[3] a_9687_8751# 0.112547f
C1073 _001_ a_5901_8751# 0.114717f
C1074 net10 _061_ 1.17544f
C1075 a_3099_9117# a_2401_8751# 0.194892f
C1076 a_1775_4399# _001_ 0.121689f
C1077 ones[9] VPWR 0.26566f
C1078 counter\[3\] VPWR 0.814878f
C1079 net5 a_3965_7663# 0.173396f
C1080 net4 net11 0.162517f
C1081 _004_ VPWR 1.86522f
C1082 _043_ net3 1.99663f
C1083 net2 net1 0.750376f
C1084 a_4491_6263# VPWR 0.181362f
C1085 _010_ counter\[8\] 0.812005f
C1086 net6 net11 0.153664f
C1087 _021_ clknet_1_1__leaf_clk 0.178906f
C1088 a_8378_9295# a_7939_9301# 0.260055f
C1089 _030_ counter\[0\] 0.107492f
C1090 a_7625_5461# counter\[5\] 0.163476f
C1091 a_4443_4949# VPWR 0.506294f
C1092 _033_ _053_ 0.352512f
C1093 counter\[8\] net11 0.198341f
C1094 a_6651_6037# clknet_1_1__leaf_clk 0.70271f
C1095 a_3965_8751# clknet_1_0__leaf_clk 0.474902f
C1096 a_8971_9269# a_8803_9295# 0.310858f
C1097 a_8767_10749# VPWR 0.432636f
C1098 _079_ _053_ 0.144407f
C1099 net7 counter\[4\] 0.882865f
C1100 _047_ _083_ 1.33016f
C1101 a_2235_8751# VPWR 0.613635f
C1102 net3 counter\[4\] 0.116331f
C1103 a_7263_7637# VPWR 0.449049f
C1104 counter\[0\] _001_ 0.18996f
C1105 ones[6] net7 0.253237f
C1106 VPWR a_9687_10927# 0.269965f
C1107 _041_ _040_ 1.14591f
C1108 a_2235_7663# _004_ 0.120991f
C1109 clk net11 0.49874f
C1110 net5 counter\[4\] 0.973692f
C1111 a_4443_4949# _006_ 0.130597f
C1112 counter\[1\] counter\[0\] 1.64337f
C1113 _002_ clknet_1_1__leaf_clk 0.191986f
C1114 net2 a_8231_4649# 0.111499f
C1115 _039_ _027_ 0.209079f
C1116 _034_ _083_ 0.153611f
C1117 a_5878_4511# VPWR 0.195622f
C1118 counter\[0\] _053_ 0.755887f
C1119 a_9411_7119# _052_ 0.139315f
C1120 a_7833_8903# _055_ 0.106268f
C1121 a_7102_6575# _018_ 0.209684f
C1122 a_8951_7663# a_9390_8029# 0.273138f
C1123 net8 net11 0.176309f
C1124 a_9687_4943# ones[7] 0.110015f
C1125 _069_ counter\[4\] 0.387961f
C1126 net7 VPWR 6.13347f
C1127 a_4319_9813# VPWR 0.389309f
C1128 net3 VPWR 3.12632f
C1129 _014_ _050_ 0.104805f
C1130 _037_ _038_ 0.109901f
C1131 _005_ _061_ 0.148549f
C1132 _070_ clknet_1_0__leaf_clk 0.599807f
C1133 _024_ counter\[5\] 0.151935f
C1134 a_9926_8181# _083_ 0.175561f
C1135 net2 a_5271_4399# 0.430847f
C1136 net5 VPWR 2.4517f
C1137 a_9648_2741# net13 0.156482f
C1138 counter\[5\] counter\[6\] 0.401086f
C1139 a_6303_4667# a_6135_4765# 0.310858f
C1140 _035_ _083_ 0.335567f
C1141 net10 net11 0.593031f
C1142 ready pulse 0.134827f
C1143 _044_ net7 0.102403f
C1144 _069_ VPWR 5.999701f
C1145 _044_ net3 0.144967f
C1146 _017_ _055_ 0.112023f
C1147 a_6411_9117# a_5713_8751# 0.191992f
C1148 a_2674_8029# VPWR 0.253282f
C1149 counter\[2\] net14 0.133648f
C1150 VPWR _045_ 0.787148f
C1151 _008_ clknet_1_1__leaf_clk 0.210761f
C1152 _007_ net12 0.515619f
C1153 a_4894_6549# a_4823_6575# 0.239923f
C1154 a_4831_7093# VPWR 0.378475f
C1155 a_7987_7828# _077_ 0.198619f
C1156 a_7711_3463# counter\[6\] 0.20796f
C1157 _005_ a_7097_4399# 0.129823f
C1158 _030_ _011_ 0.108856f
C1159 a_10199_3285# VPWR 0.369039f
C1160 a_6814_8207# a_6375_8213# 0.260055f
C1161 _037_ a_2509_4663# 0.214381f
C1162 _014_ net12 0.350809f
C1163 a_7090_6031# VPWR 0.255868f
C1164 _040_ _053_ 0.134874f
C1165 counter\[1\] net13 0.391575f
C1166 a_9963_10383# ones[10] 0.111194f
C1167 a_6189_6825# VPWR 0.1903f
C1168 net4 _049_ 0.145261f
C1169 _072_ _042_ 0.149428f
C1170 a_2674_8029# a_2235_7663# 0.273138f
C1171 _083_ net12 0.272125f
C1172 a_9551_9527# _086_ 0.196759f
C1173 a_2409_5263# counter\[10\] 0.173455f
C1174 a_2431_5487# VPWR 0.180149f
C1175 _047_ _051_ 0.281094f
C1176 net6 a_8268_2741# 0.122657f
C1177 clknet_1_1__leaf_clk counter\[2\] 0.127194f
C1178 _037_ _021_ 0.172905f
C1179 a_7987_7351# net6 0.108608f
C1180 _065_ VPWR 1.2006f
C1181 _023_ _045_ 0.1269f
C1182 _064_ counter\[5\] 0.221545f
C1183 _055_ _050_ 0.199126f
C1184 _084_ _004_ 1.11974f
C1185 a_9739_6005# _028_ 0.12491f
C1186 a_9963_10383# VPWR 0.260504f
C1187 a_4687_6549# clknet_0_clk 0.101639f
C1188 a_9411_7119# _050_ 0.109782f
C1189 _009_ net6 0.126615f
C1190 a_4403_6549# VPWR 0.171892f
C1191 _054_ VPWR 0.739884f
C1192 counter\[1\] counter\[3\] 0.470344f
C1193 _013_ _052_ 0.230849f
C1194 a_5475_4917# a_5307_4943# 0.310858f
C1195 clknet_1_0__leaf_clk _086_ 1.01249f
C1196 a_10134_10927# counter\[8\] 0.184047f
C1197 _027_ VPWR 1.86707f
C1198 _069_ _025_ 0.115762f
C1199 net2 _040_ 0.456288f
C1200 a_4801_10973# _027_ 0.123111f
C1201 _069_ _041_ 0.480687f
C1202 _078_ VPWR 1.78731f
C1203 a_4491_6263# _053_ 0.181294f
C1204 a_9926_8181# net14 0.214732f
C1205 a_4981_6263# _036_ 0.101875f
C1206 net9 _077_ 0.88188f
C1207 net2 net13 0.81239f
C1208 _014_ a_3799_7125# 0.427292f
C1209 a_5547_8751# counter\[8\] 0.106769f
C1210 counter\[7\] a_3867_9813# 0.12818f
C1211 _051_ _050_ 0.661737f
C1212 a_2787_4949# a_2953_4949# 0.960876f
C1213 net4 _036_ 0.858449f
C1214 a_3965_8751# a_3799_8751# 0.961627f
C1215 a_4831_9019# a_4663_9117# 0.310858f
C1216 _035_ _051_ 0.297172f
C1217 _044_ _027_ 0.923831f
C1218 _071_ counter\[8\] 0.294774f
C1219 a_1573_9839# VPWR 0.358186f
C1220 _044_ _078_ 3.40291f
C1221 _063_ _062_ 1.80289f
C1222 a_9390_8029# VPWR 0.253921f
C1223 _043_ _075_ 0.236947f
C1224 clknet_1_0__leaf_clk a_4326_10113# 0.456134f
C1225 _043_ _058_ 0.137772f
C1226 net2 counter\[3\] 0.104721f
C1227 a_2842_8863# VPWR 0.178412f
C1228 a_4589_3829# VPWR 0.206652f
C1229 a_3799_7663# _000_ 0.122534f
C1230 a_4406_8863# a_4238_9117# 0.239923f
C1231 _021_ _086_ 0.305801f
C1232 a_9305_6575# _018_ 0.114994f
C1233 counter\[1\] net3 0.698949f
C1234 ones[7] VPWR 0.37058f
C1235 clknet_1_1__leaf_clk _050_ 0.157826f
C1236 _084_ net5 0.142528f
C1237 _024_ _026_ 0.105485f
C1238 _070_ counter\[9\] 0.110956f
C1239 net7 _053_ 0.234921f
C1240 _027_ a_1761_2999# 0.100598f
C1241 net3 _053_ 0.263248f
C1242 _085_ _022_ 0.130688f
C1243 _061_ net11 0.277724f
C1244 _066_ _035_ 0.785244f
C1245 net5 counter\[1\] 0.242765f
C1246 _037_ counter\[7\] 0.520583f
C1247 net12 net14 0.360111f
C1248 net1 net14 1.36538f
C1249 a_5496_9269# _042_ 0.115867f
C1250 a_7939_9301# clknet_1_1__leaf_clk 0.22857f
C1251 net5 _053_ 0.219753f
C1252 _069_ _001_ 0.782639f
C1253 a_6511_5461# counter\[0\] 0.226488f
C1254 _025_ _027_ 0.337557f
C1255 clknet_1_1__leaf_clk a_8367_7337# 0.672881f
C1256 net12 _051_ 0.18139f
C1257 a_9247_6005# net4 0.148333f
C1258 _026_ _086_ 0.16073f
C1259 a_4455_9839# VPWR 0.174858f
C1260 _035_ _028_ 0.195238f
C1261 a_4443_4949# a_5050_4917# 0.136009f
C1262 _069_ counter\[1\] 0.308236f
C1263 _052_ a_8374_7241# 0.36233f
C1264 a_9815_6941# a_9983_6843# 0.310858f
C1265 _076_ a_8374_7241# 0.114034f
C1266 _069_ _053_ 0.406937f
C1267 a_2302_5761# counter\[9\] 0.187019f
C1268 _071_ net10 0.107447f
C1269 a_8215_6037# net7 0.436809f
C1270 _002_ net9 0.104906f
C1271 _075_ VPWR 2.80706f
C1272 _058_ VPWR 1.97125f
C1273 a_4135_4373# _061_ 0.123346f
C1274 _016_ a_5271_8751# 0.109137f
C1275 _036_ net10 0.288393f
C1276 net2 net3 0.652313f
C1277 net4 counter\[5\] 0.663311f
C1278 a_8231_4649# net14 0.116858f
C1279 net12 clknet_1_1__leaf_clk 0.125777f
C1280 net1 clknet_1_1__leaf_clk 0.142367f
C1281 _063_ counter\[4\] 0.197836f
C1282 _073_ counter\[3\] 0.250962f
C1283 _080_ _035_ 1.91257f
C1284 _013_ a_8367_7337# 0.102104f
C1285 net6 counter\[5\] 0.167155f
C1286 net2 net5 0.165127f
C1287 _067_ VPWR 0.714476f
C1288 counter\[5\] counter\[8\] 0.108937f
C1289 _020_ _061_ 0.692663f
C1290 a_2787_4949# _079_ 0.100522f
C1291 _024_ counter\[7\] 0.89735f
C1292 counter\[0\] _055_ 0.159928f
C1293 _001_ _065_ 0.261142f
C1294 a_9011_3285# _086_ 0.172852f
C1295 _024_ counter\[9\] 0.783525f
C1296 _016_ _017_ 0.102183f
C1297 net12 _028_ 0.422524f
C1298 _033_ _051_ 0.245434f
C1299 net1 _028_ 0.423534f
C1300 a_9011_3285# _031_ 0.190477f
C1301 _012_ VPWR 0.497404f
C1302 _005_ a_6909_4399# 0.199131f
C1303 _083_ net13 0.115071f
C1304 a_7515_6031# VPWR 0.17179f
C1305 counter\[7\] counter\[6\] 2.13747f
C1306 a_4621_10383# VPWR 0.248927f
C1307 _056_ _009_ 0.270068f
C1308 _018_ _055_ 0.774496f
C1309 _007_ counter\[3\] 0.105323f
C1310 a_3421_3855# VPWR 0.166242f
C1311 a_4798_5737# counter\[2\] 0.111141f
C1312 net9 a_9011_3285# 0.197668f
C1313 _053_ _065_ 1.04867f
C1314 _008_ _031_ 0.331391f
C1315 clk counter\[5\] 0.1003f
C1316 _023_ _075_ 0.475071f
C1317 _058_ _023_ 0.821573f
C1318 counter\[7\] _086_ 0.334228f
C1319 _063_ VPWR 1.99942f
C1320 _013_ a_8921_7497# 0.114667f
C1321 _046_ _036_ 0.128095f
C1322 a_6982_8181# a_6814_8207# 0.239923f
C1323 counter\[7\] _031_ 0.105153f
C1324 counter\[10\] VPWR 2.34698f
C1325 net9 _008_ 0.412042f
C1326 clknet_0_clk counter\[4\] 0.308481f
C1327 a_8381_6037# VPWR 0.276595f
C1328 _084_ _078_ 0.540056f
C1329 counter\[9\] _086_ 0.63635f
C1330 _001_ _078_ 1.1285f
C1331 _076_ counter\[6\] 0.666412f
C1332 _054_ _053_ 0.124984f
C1333 net9 counter\[7\] 0.346546f
C1334 a_4351_5737# VPWR 0.32168f
C1335 a_3267_9019# VPWR 0.399921f
C1336 _024_ counter\[2\] 0.119134f
C1337 _072_ VPWR 3.4647f
C1338 a_7258_6005# a_6651_6037# 0.135468f
C1339 counter\[1\] _078_ 0.184242f
C1340 _076_ _086_ 0.182535f
C1341 _080_ net1 0.296532f
C1342 a_2011_5461# VPWR 0.186474f
C1343 a_4406_7775# a_3799_7663# 0.136009f
C1344 _083_ counter\[3\] 1.17069f
C1345 counter\[6\] counter\[2\] 0.782721f
C1346 a_4687_6549# VPWR 0.584529f
C1347 net9 _076_ 0.254729f
C1348 _042_ VPWR 0.684196f
C1349 counter\[2\] _086_ 0.198305f
C1350 a_5271_4399# clknet_1_1__leaf_clk 0.293108f
C1351 net9 a_9739_6005# 0.157378f
C1352 a_9117_6575# a_9558_6687# 0.124967f
C1353 a_7829_4949# VPWR 0.276911f
C1354 a_2014_9951# a_1846_10205# 0.239923f
C1355 clknet_0_clk VPWR 3.20387f
C1356 a_8953_2473# VPWR 0.269352f
C1357 clknet_1_0__leaf_clk a_2401_8751# 0.377366f
C1358 net10 counter\[5\] 0.2466f
C1359 _024_ _017_ 0.333466f
C1360 a_4120_3291# _024_ 0.102104f
C1361 _059_ counter\[0\] 1.17691f
C1362 a_2409_5263# VPWR 0.1733f
C1363 _047_ _024_ 0.166514f
C1364 clknet_1_0__leaf_clk counter\[8\] 0.360748f
C1365 _043_ _039_ 0.131887f
C1366 _029_ _056_ 0.614343f
C1367 _085_ _064_ 0.416195f
C1368 _040_ _055_ 0.456059f
C1369 counter\[0\] clknet_1_1__leaf_clk 0.673232f
C1370 _069_ _073_ 0.205315f
C1371 a_2787_4949# a_3226_4943# 0.260055f
C1372 a_2953_4949# a_3394_4917# 0.110715f
C1373 _015_ counter\[2\] 0.509654f
C1374 a_8367_7337# a_8374_7241# 0.960615f
C1375 a_3137_4765# VPWR 0.335428f
C1376 net8 a_9551_9527# 0.168329f
C1377 _074_ counter\[9\] 0.220525f
C1378 a_9687_4943# VPWR 0.258264f
C1379 _081_ net1 0.127201f
C1380 VPWR a_7607_4765# 0.184612f
C1381 a_4120_3291# _031_ 0.119534f
C1382 _047_ _086_ 0.212279f
C1383 clknet_1_1__leaf_clk _018_ 0.739046f
C1384 a_9815_8029# VPWR 0.193764f
C1385 a_8270_4917# a_7829_4949# 0.110715f
C1386 _047_ _031_ 0.211452f
C1387 a_3847_3463# _024_ 0.115316f
C1388 a_4798_5737# _050_ 0.195074f
C1389 _034_ a_3851_6005# 0.107169f
C1390 _030_ _058_ 0.969056f
C1391 a_5607_10089# VPWR 0.190299f
C1392 a_8355_4074# VPWR 0.234599f
C1393 a_8951_7663# VPWR 0.620401f
C1394 _069_ _007_ 0.470417f
C1395 a_4234_9417# _042_ 0.105386f
C1396 _083_ net3 1.31226f
C1397 _034_ _086_ 0.47328f
C1398 VPWR rst 0.305657f
C1399 _021_ net4 0.261618f
C1400 a_2143_7232# VPWR 0.240845f
C1401 net13 net14 0.491806f
C1402 net5 _083_ 0.679661f
C1403 _024_ _035_ 0.2581f
C1404 ones[7] ready 0.176502f
C1405 a_5713_8751# a_6154_8863# 0.110715f
C1406 counter\[1\] _075_ 0.10942f
C1407 _080_ counter\[0\] 0.354252f
C1408 _058_ counter\[1\] 0.185964f
C1409 a_3847_6727# _061_ 0.210887f
C1410 _039_ VPWR 4.25447f
C1411 a_6135_4765# a_5437_4399# 0.192261f
C1412 _062_ VPWR 1.18935f
C1413 _069_ _083_ 0.195862f
C1414 _075_ _053_ 0.151201f
C1415 _058_ _053_ 0.242609f
C1416 a_3965_8751# a_4406_8863# 0.110715f
C1417 a_9735_5639# _085_ 0.120815f
C1418 a_5496_9269# VPWR 0.208821f
C1419 _059_ net13 0.338038f
C1420 _010_ _049_ 0.52719f
C1421 _040_ clknet_1_1__leaf_clk 0.265958f
C1422 a_3203_7351# VPWR 0.198332f
C1423 a_3651_4943# a_2953_4949# 0.192261f
C1424 a_3965_7125# a_3799_7125# 0.961627f
C1425 _045_ a_2419_2767# 0.113506f
C1426 a_7939_9301# _086_ 0.108765f
C1427 a_4601_5737# a_4798_5737# 0.149348f
C1428 _084_ _012_ 0.634441f
C1429 _067_ _053_ 0.165686f
C1430 _012_ _001_ 0.483168f
C1431 _044_ _039_ 0.294581f
C1432 _015_ _050_ 0.694842f
C1433 a_3867_9813# a_4035_9813# 0.310858f
C1434 _067_ a_5823_7119# 0.189319f
C1435 _060_ a_6375_2767# 0.194319f
C1436 _024_ net1 0.223354f
C1437 VPWR a_7531_2741# 0.186622f
C1438 a_3965_7663# VPWR 0.277325f
C1439 _012_ _053_ 0.103711f
C1440 a_7616_7351# VPWR 0.16044f
C1441 counter\[1\] _063_ 0.153995f
C1442 net3 _055_ 0.113578f
C1443 _072_ _001_ 0.229896f
C1444 net1 counter\[6\] 0.76912f
C1445 a_9503_8207# net5 0.195295f
C1446 _043_ VPWR 1.59127f
C1447 a_4351_5737# counter\[1\] 0.136251f
C1448 _021_ net10 1.5876f
C1449 net12 _086_ 0.159731f
C1450 ones[0] net13 0.169258f
C1451 net1 _086_ 0.193712f
C1452 net12 _031_ 0.451082f
C1453 VPWR a_6743_4399# 0.436963f
C1454 net1 _031_ 0.280414f
C1455 _035_ _074_ 0.435238f
C1456 _072_ _053_ 0.196433f
C1457 _071_ net11 0.220754f
C1458 a_2787_6031# _024_ 0.134565f
C1459 _016_ counter\[0\] 0.126937f
C1460 a_5433_7637# net1 0.145917f
C1461 net7 net14 0.433924f
C1462 _025_ _039_ 2.13004f
C1463 _027_ _083_ 0.265955f
C1464 _036_ net11 0.102094f
C1465 a_3965_7125# a_4406_7093# 0.110715f
C1466 net3 net14 0.398434f
C1467 _020_ _049_ 0.607312f
C1468 counter\[5\] _061_ 0.36662f
C1469 a_7102_6575# clknet_0_clk 0.327485f
C1470 a_8231_4649# _024_ 0.152804f
C1471 ones[2] net1 0.193638f
C1472 counter\[4\] VPWR 4.24859f
C1473 net7 _051_ 1.34574f
C1474 _053_ _042_ 0.211206f
C1475 ones[8] a_9687_8751# 0.110363f
C1476 a_7829_4949# _053_ 0.371076f
C1477 a_6979_10901# VPWR 0.307879f
C1478 counter\[7\] counter\[8\] 0.942849f
C1479 ones[10] VPWR 0.154188f
C1480 net5 net14 0.216405f
C1481 ones[6] VPWR 0.385576f
C1482 a_3819_4917# a_3651_4943# 0.310858f
C1483 a_8215_6037# a_8381_6037# 0.961627f
C1484 counter\[9\] counter\[8\] 0.388388f
C1485 _024_ _033_ 0.122641f
C1486 _052_ net6 0.297664f
C1487 a_6060_6549# VPWR 0.213251f
C1488 net6 _076_ 0.231801f
C1489 _076_ counter\[8\] 0.113702f
C1490 a_9558_6687# a_9390_6941# 0.239923f
C1491 _033_ counter\[6\] 0.469288f
C1492 _003_ a_2401_8751# 0.198156f
C1493 _021_ _046_ 0.199238f
C1494 net8 a_9011_3285# 0.156282f
C1495 _069_ _051_ 0.743064f
C1496 _009_ a_4227_9513# 0.134448f
C1497 a_9079_6031# a_8381_6037# 0.192261f
C1498 net7 clknet_1_1__leaf_clk 0.612806f
C1499 a_4801_10973# VPWR 0.175247f
C1500 _074_ net1 0.133475f
C1501 net3 clknet_1_1__leaf_clk 0.283214f
C1502 counter\[2\] counter\[8\] 0.685145f
C1503 clk _076_ 0.291033f
C1504 a_3394_4917# a_3226_4943# 0.239923f
C1505 _070_ _040_ 0.238337f
C1506 _024_ counter\[0\] 0.108746f
C1507 a_8367_7337# a_8503_7497# 0.136009f
C1508 a_5043_4564# VPWR 0.190083f
C1509 a_9411_8751# net7 0.221455f
C1510 net5 clknet_1_1__leaf_clk 0.170705f
C1511 VPWR a_10239_4399# 0.216414f
C1512 _021_ _056_ 0.125897f
C1513 _054_ a_2879_8207# 0.190426f
C1514 _006_ VPWR 0.330292f
C1515 _044_ VPWR 2.85077f
C1516 a_2143_7232# _053_ 0.168735f
C1517 _037_ _040_ 0.321915f
C1518 net10 _008_ 1.02271f
C1519 a_8270_4917# VPWR 0.176131f
C1520 a_2235_7663# VPWR 0.65145f
C1521 net10 _085_ 0.124364f
C1522 net5 _028_ 0.832261f
C1523 net8 a_9739_6005# 0.153151f
C1524 a_8654_6031# VPWR 0.242357f
C1525 net10 counter\[7\] 0.101175f
C1526 a_7663_4949# a_7829_4949# 0.961627f
C1527 a_2302_5761# a_2295_5461# 0.973502f
C1528 _010_ counter\[5\] 0.110552f
C1529 ones[0] net3 0.208275f
C1530 _013_ net7 0.705811f
C1531 a_5271_4399# a_5437_4399# 0.961627f
C1532 _023_ VPWR 3.44101f
C1533 _039_ _053_ 0.477692f
C1534 _018_ _086_ 0.110952f
C1535 counter\[5\] net11 0.201202f
C1536 net9 pulse 0.392665f
C1537 _025_ ones[10] 0.144734f
C1538 _011_ _016_ 0.153599f
C1539 net3 _060_ 1.19532f
C1540 a_4238_8029# VPWR 0.237894f
C1541 a_4234_9417# VPWR 0.304546f
C1542 _083_ _075_ 0.163688f
C1543 _080_ net3 0.475574f
C1544 a_1761_2999# VPWR 0.194512f
C1545 a_6154_8863# a_5986_9117# 0.239923f
C1546 _034_ counter\[8\] 0.242112f
C1547 clknet_1_0__leaf_clk a_3799_7663# 0.228232f
C1548 a_9735_5639# net1 0.194733f
C1549 a_8091_10615# VPWR 0.217317f
C1550 _079_ _064_ 1.20609f
C1551 a_4609_4949# a_5307_4943# 0.194215f
C1552 _044_ _023_ 0.487411f
C1553 _025_ VPWR 2.83838f
C1554 clknet_1_0__leaf_clk _000_ 0.674307f
C1555 _041_ VPWR 0.44777f
C1556 net4 _035_ 0.185535f
C1557 net8 _047_ 0.233241f
C1558 _048_ _050_ 0.36959f
C1559 a_6743_4399# a_7350_4511# 0.136009f
C1560 _083_ _067_ 0.436448f
C1561 a_4035_9813# a_4326_10113# 0.192261f
C1562 _048_ _035_ 0.318546f
C1563 _024_ _040_ 0.594233f
C1564 a_4238_7119# a_3799_7125# 0.260055f
C1565 net2 _039_ 0.216797f
C1566 counter\[0\] _068_ 0.140058f
C1567 _035_ counter\[8\] 0.107445f
C1568 _021_ _061_ 1.34574f
C1569 a_5731_3311# VPWR 0.224782f
C1570 _043_ _053_ 0.400131f
C1571 _068_ _018_ 0.153262f
C1572 _020_ counter\[5\] 0.531736f
C1573 VPWR a_9648_2741# 0.21022f
C1574 _063_ a_3479_10004# 0.214865f
C1575 ones[8] net13 0.885732f
C1576 a_4227_9513# a_4434_9572# 0.273138f
C1577 a_8083_7351# VPWR 0.178379f
C1578 clknet_1_1__leaf_clk _078_ 0.102972f
C1579 _019_ a_2007_7828# 0.108595f
C1580 _010_ clknet_1_0__leaf_clk 0.687869f
C1581 clknet_1_0__leaf_clk net11 0.163469f
C1582 a_5503_11092# VPWR 0.248794f
C1583 _082_ counter\[0\] 0.134668f
C1584 a_2401_7663# a_3099_8029# 0.194892f
C1585 a_7407_8181# a_7239_8207# 0.310858f
C1586 _077_ net11 1.06665f
C1587 _030_ VPWR 0.559897f
C1588 net8 _050_ 0.26514f
C1589 _024_ counter\[3\] 0.192447f
C1590 _056_ _052_ 0.324262f
C1591 _053_ counter\[4\] 0.436151f
C1592 _022_ net7 0.321621f
C1593 VPWR a_7350_4511# 0.19494f
C1594 _037_ net7 0.128422f
C1595 net8 _035_ 0.13832f
C1596 net4 net1 0.775071f
C1597 _014_ clknet_0_clk 0.115783f
C1598 a_6099_10089# _004_ 0.101082f
C1599 net12 net6 0.705267f
C1600 net6 net1 0.17515f
C1601 a_3847_3463# _032_ 0.20232f
C1602 a_2401_7663# a_2842_7775# 0.110174f
C1603 a_9861_5737# VPWR 0.202725f
C1604 _030_ a_5043_4564# 0.191318f
C1605 a_2143_7232# _073_ 0.210182f
C1606 _069_ _070_ 0.359237f
C1607 a_4406_7093# a_4238_7119# 0.239923f
C1608 net12 counter\[8\] 0.20143f
C1609 _084_ VPWR 2.73277f
C1610 _013_ _027_ 0.167867f
C1611 _001_ VPWR 1.24989f
C1612 a_10199_2197# rst 0.250422f
C1613 _004_ _086_ 0.385541f
C1614 a_7102_6575# VPWR 1.28968f
C1615 VPWR a_2439_10107# 0.471319f
C1616 a_7515_6031# a_6817_6037# 0.191064f
C1617 _047_ _046_ 0.146843f
C1618 net10 _050_ 0.144837f
C1619 a_4694_6849# _017_ 0.188635f
C1620 counter\[1\] VPWR 2.14401f
C1621 net2 a_6743_4399# 0.442672f
C1622 a_3847_9527# VPWR 0.394436f
C1623 _038_ _020_ 1.12944f
C1624 _069_ _016_ 0.465542f
C1625 a_4663_8029# a_3965_7663# 0.192261f
C1626 _053_ VPWR 7.66588f
C1627 clk net12 0.460451f
C1628 a_5823_7119# VPWR 0.238677f
C1629 ones[3] VPWR 0.422382f
C1630 _084_ _044_ 0.137777f
C1631 _044_ _001_ 0.37197f
C1632 a_2409_4445# VPWR 0.178195f
C1633 a_7263_7637# _086_ 0.154026f
C1634 _085_ _061_ 0.107758f
C1635 _011_ _074_ 0.108858f
C1636 net8 net1 0.107704f
C1637 a_4694_6849# a_4823_6575# 0.112272f
C1638 a_4687_6549# a_4894_6549# 0.271965f
C1639 _024_ net7 0.146913f
C1640 counter\[7\] _061_ 0.552061f
C1641 a_9117_6575# a_8951_6575# 0.967319f
C1642 _044_ _053_ 1.8136f
C1643 ready VPWR 0.205435f
C1644 a_3137_4765# a_2971_4399# 0.124682f
C1645 a_8574_7396# a_8503_7497# 0.239923f
C1646 clknet_1_0__leaf_clk a_4227_9513# 0.229782f
C1647 a_3851_6005# net7 0.177396f
C1648 _070_ _065_ 0.166195f
C1649 a_8215_6037# VPWR 0.429228f
C1650 net7 counter\[6\] 0.38915f
C1651 _076_ _061_ 0.646444f
C1652 _004_ a_6324_10029# 0.146368f
C1653 net2 VPWR 4.88291f
C1654 net7 _086_ 1.68994f
C1655 _023_ _053_ 1.96862f
C1656 net10 net12 0.832341f
C1657 net3 _086_ 0.369147f
C1658 net10 net1 0.129353f
C1659 net5 counter\[6\] 0.114068f
C1660 _011_ _082_ 0.122591f
C1661 a_8695_4917# VPWR 0.388551f
C1662 ready a_10239_4399# 0.11283f
C1663 _069_ _024_ 1.19048f
C1664 net9 net7 0.114756f
C1665 a_9079_6031# VPWR 0.169797f
C1666 net9 net3 0.23519f
C1667 net3 a_5433_7637# 0.115498f
C1668 net5 _086_ 1.17506f
C1669 VPWR a_10239_8751# 0.274041f
C1670 a_2295_5461# a_2502_5461# 0.273138f
C1671 a_2302_5761# a_2431_5487# 0.117154f
C1672 a_5437_4399# a_5878_4511# 0.110715f
C1673 a_5271_4399# a_5710_4765# 0.260055f
C1674 _038_ _049_ 0.427615f
C1675 _039_ a_2419_2767# 0.131238f
C1676 a_7663_4949# VPWR 0.414564f
C1677 _069_ counter\[6\] 0.292105f
C1678 a_5050_4917# VPWR 0.174439f
C1679 _035_ _057_ 0.289857f
C1680 counter\[0\] counter\[8\] 0.488018f
C1681 net5 a_5433_7637# 0.213066f
C1682 a_4663_8029# VPWR 0.172668f
C1683 a_5018_5461# _050_ 0.136664f
C1684 a_4363_9673# VPWR 0.182441f
C1685 a_8654_6031# a_8215_6037# 0.260055f
C1686 a_3847_6727# counter\[5\] 0.166922f
C1687 a_1673_10973# VPWR 0.179608f
C1688 clknet_1_0__leaf_clk _049_ 0.288759f
C1689 _018_ counter\[8\] 0.120635f
C1690 a_2302_5761# _027_ 0.101568f
C1691 _069_ net9 0.402552f
C1692 a_8378_9295# VPWR 0.260183f
C1693 _058_ _060_ 0.109776f
C1694 a_4326_10113# a_4319_9813# 0.961627f
C1695 _046_ net1 0.43894f
C1696 a_8546_9269# a_8105_9301# 0.110715f
C1697 _069_ _015_ 0.250197f
C1698 a_8270_4917# a_7663_4949# 0.136009f
C1699 _074_ net7 0.216521f
C1700 clknet_1_0__leaf_clk _009_ 0.28314f
C1701 net7 _064_ 0.221084f
C1702 _012_ a_4153_8751# 0.114652f
C1703 counter\[7\] net11 0.128533f
C1704 _010_ counter\[9\] 0.153223f
C1705 net8 counter\[0\] 0.389654f
C1706 a_2776_7119# _026_ 0.164723f
C1707 _034_ _061_ 0.150437f
C1708 _073_ VPWR 1.62765f
C1709 a_8075_3285# VPWR 0.232925f
C1710 a_6979_10901# _007_ 0.10607f
C1711 net8 pulse 0.20348f
C1712 a_3137_4765# _051_ 0.191345f
C1713 a_4687_6549# clknet_1_1__leaf_clk 0.316547f
C1714 counter\[6\] _065_ 0.193763f
C1715 _024_ _054_ 0.258083f
C1716 _043_ a_2419_2767# 0.138082f
C1717 a_10199_2197# VPWR 0.375761f
C1718 a_6375_8213# VPWR 0.480025f
C1719 _046_ a_2787_6031# 0.1394f
C1720 a_8123_5487# net6 0.141239f
C1721 _014_ counter\[4\] 0.154626f
C1722 clknet_1_0__leaf_clk a_5547_8751# 0.221375f
C1723 _024_ _027_ 1.54154f
C1724 _062_ _055_ 0.718567f
C1725 a_4234_9417# a_4363_9673# 0.110715f
C1726 net4 _040_ 0.393617f
C1727 _069_ _074_ 0.102216f
C1728 _069_ _068_ 0.130839f
C1729 a_2051_4943# counter\[7\] 0.112207f
C1730 a_10103_9514# VPWR 0.229526f
C1731 net10 counter\[0\] 0.152185f
C1732 a_9117_7663# a_9558_7775# 0.124967f
C1733 net6 _040_ 0.218562f
C1734 net4 net13 0.972738f
C1735 _061_ _050_ 0.200878f
C1736 _007_ VPWR 0.518287f
C1737 _054_ _086_ 0.1537f
C1738 _029_ _038_ 0.560511f
C1739 counter\[2\] net11 0.124497f
C1740 _084_ _053_ 0.135299f
C1741 _012_ a_3965_8751# 0.180738f
C1742 a_6411_9117# VPWR 0.168006f
C1743 _027_ _086_ 0.87618f
C1744 counter\[8\] net13 0.156101f
C1745 _086_ _078_ 0.139199f
C1746 _014_ VPWR 1.65571f
C1747 _027_ net9 0.113405f
C1748 a_2842_7775# a_2674_8029# 0.239923f
C1749 a_10103_9991# VPWR 0.238437f
C1750 _020_ counter\[7\] 0.162194f
C1751 a_9735_5639# net3 0.110955f
C1752 VPWR a_3479_10004# 0.26833f
C1753 _083_ VPWR 3.17235f
C1754 _082_ _045_ 0.420057f
C1755 a_8951_7663# clknet_1_1__leaf_clk 0.218176f
C1756 a_4238_9117# VPWR 0.240909f
C1757 a_5241_6575# _017_ 0.121794f
C1758 a_8951_6575# _018_ 0.137728f
C1759 a_1775_4399# _057_ 0.190667f
C1760 a_4443_4949# a_4609_4949# 0.973227f
C1761 a_4135_4373# counter\[2\] 0.159185f
C1762 _056_ _033_ 0.857459f
C1763 _020_ _052_ 0.151199f
C1764 VPWR a_2419_2767# 0.639838f
C1765 a_9735_5639# net5 0.122703f
C1766 a_6511_5461# VPWR 0.203406f
C1767 a_2971_4399# VPWR 0.19221f
C1768 net12 _061_ 0.787649f
C1769 net2 counter\[1\] 0.134383f
C1770 _021_ _036_ 0.100282f
C1771 _027_ _068_ 0.310501f
C1772 a_9390_6941# a_8951_6575# 0.260364f
C1773 a_2235_8751# a_2401_8751# 0.961428f
C1774 a_7258_6005# a_7090_6031# 0.239923f
C1775 a_6303_4667# VPWR 0.374997f
C1776 a_7263_7637# net6 0.15825f
C1777 _044_ a_2419_2767# 0.159072f
C1778 net10 _040_ 0.308741f
C1779 _025_ a_10103_9514# 0.190836f
C1780 _056_ counter\[0\] 0.295889f
C1781 _010_ a_3593_8181# 0.172322f
C1782 _023_ _083_ 0.413587f
C1783 a_5018_5461# counter\[0\] 0.160435f
C1784 a_4894_6549# VPWR 0.253369f
C1785 ones[7] ones[2] 0.206144f
C1786 a_6817_6037# VPWR 0.292675f
C1787 a_4807_3855# VPWR 0.222624f
C1788 a_2734_6575# net11 0.105614f
C1789 _058_ _024_ 0.431245f
C1790 _035_ net11 0.718948f
C1791 net4 net7 0.138281f
C1792 a_9117_6575# net11 0.147779f
C1793 _077_ counter\[5\] 0.511495f
C1794 ones[1] VPWR 0.343002f
C1795 net4 net3 0.978794f
C1796 counter\[7\] _049_ 0.601021f
C1797 net2 ready 0.24238f
C1798 a_9503_8207# VPWR 0.216403f
C1799 _075_ counter\[6\] 0.102795f
C1800 net7 net6 0.128756f
C1801 a_2879_8207# VPWR 0.27095f
C1802 counter\[9\] _049_ 0.102048f
C1803 net3 net6 0.708983f
C1804 a_2502_5461# a_2431_5487# 0.239923f
C1805 _055_ VPWR 1.17426f
C1806 _043_ _059_ 1.43435f
C1807 a_5878_4511# a_5710_4765# 0.239923f
C1808 counter\[4\] _051_ 0.278002f
C1809 _049_ _052_ 1.61727f
C1810 a_9411_7119# VPWR 0.590119f
C1811 _024_ _067_ 0.402798f
C1812 a_5475_4917# VPWR 0.391553f
C1813 _033_ _061_ 0.111237f
C1814 a_5363_6031# VPWR 0.189968f
C1815 _049_ _076_ 0.107086f
C1816 net5 net6 1.61745f
C1817 a_2302_5761# a_2011_5461# 0.193199f
C1818 _016_ clknet_0_clk 0.690011f
C1819 a_4781_9673# _009_ 0.114852f
C1820 _079_ _061_ 0.140915f
C1821 a_2787_4949# VPWR 0.436972f
C1822 clknet_1_1__leaf_clk a_6743_4399# 0.302405f
C1823 a_3476_7351# a_3203_7351# 0.167615f
C1824 clk net7 0.193178f
C1825 _069_ _048_ 0.486354f
C1826 net4 _045_ 0.340465f
C1827 a_8803_9295# VPWR 0.18616f
C1828 a_4326_10113# a_4455_9839# 0.110715f
C1829 a_4319_9813# a_4526_9813# 0.260055f
C1830 VPWR net14 1.31648f
C1831 _069_ counter\[8\] 3.5362f
C1832 a_4307_6727# a_4403_6549# 0.310858f
C1833 _024_ counter\[10\] 1.27643f
C1834 net12 net11 0.884528f
C1835 net1 net11 0.35774f
C1836 VPWR _051_ 1.34687f
C1837 _057_ _040_ 0.108088f
C1838 clknet_1_1__leaf_clk counter\[4\] 0.457135f
C1839 net8 net7 0.426708f
C1840 _071_ counter\[7\] 0.297454f
C1841 _066_ counter\[4\] 0.295609f
C1842 _019_ a_1761_9839# 0.137291f
C1843 a_8293_9295# _022_ 0.12468f
C1844 _071_ a_7108_5737# 0.113934f
C1845 ones[10] ones[4] 0.17677f
C1846 a_10239_10383# ones[10] 0.117773f
C1847 _018_ _061_ 0.59968f
C1848 _022_ a_8355_4074# 0.122157f
C1849 counter\[10\] _086_ 0.386722f
C1850 _068_ _075_ 0.16533f
C1851 _059_ VPWR 0.631068f
C1852 _043_ _060_ 0.331736f
C1853 _011_ a_3141_4943# 0.124835f
C1854 _024_ _042_ 0.305754f
C1855 _075_ _064_ 1.01314f
C1856 _058_ _068_ 0.431396f
C1857 a_8727_8181# _078_ 0.120428f
C1858 a_2014_9951# a_1407_9839# 0.141453f
C1859 _029_ _085_ 0.238795f
C1860 net10 net7 0.228874f
C1861 _072_ _086_ 0.111479f
C1862 _070_ _039_ 0.526819f
C1863 net10 net3 0.926999f
C1864 a_9983_7931# net13 0.156988f
C1865 clknet_1_1__leaf_clk VPWR 5.22238f
C1866 a_2674_9117# a_2235_8751# 0.273138f
C1867 _032_ net3 0.122614f
C1868 _048_ _065_ 0.237184f
C1869 net4 a_9963_10383# 0.224573f
C1870 a_6541_8213# _008_ 0.261259f
C1871 ones[4] VPWR 0.409295f
C1872 _066_ VPWR 0.26362f
C1873 a_10239_10383# VPWR 0.216102f
C1874 a_10103_9991# _053_ 0.167446f
C1875 net5 net10 0.173636f
C1876 _042_ _086_ 0.164792f
C1877 _074_ _067_ 1.16392f
C1878 a_6982_8181# VPWR 0.193717f
C1879 counter\[1\] _083_ 0.285668f
C1880 a_7683_6005# net7 0.137277f
C1881 _065_ counter\[8\] 0.312238f
C1882 net2 a_10199_2197# 0.177245f
C1883 a_9411_8751# VPWR 0.231708f
C1884 _083_ _053_ 1.84672f
C1885 a_4491_6263# _056_ 0.199516f
C1886 VPWR _028_ 0.831401f
C1887 clknet_0_clk a_5433_7637# 1.63724f
C1888 _029_ counter\[2\] 0.163705f
C1889 _049_ _050_ 2.45675f
C1890 a_6511_5461# _053_ 0.128072f
C1891 ones[0] VPWR 0.181336f
C1892 a_4153_7119# _015_ 0.12469f
C1893 a_4831_7093# a_4663_7119# 0.310858f
C1894 _078_ counter\[8\] 0.171261f
C1895 _032_ _045_ 0.71586f
C1896 _035_ _049_ 0.237705f
C1897 a_4663_9117# VPWR 0.171738f
C1898 _064_ _063_ 0.121208f
C1899 _013_ VPWR 0.607678f
C1900 _046_ net7 1.25932f
C1901 _074_ counter\[10\] 0.172708f
C1902 _040_ _061_ 0.406155f
C1903 a_9558_7775# a_9390_8029# 0.239923f
C1904 _010_ counter\[0\] 0.256011f
C1905 a_3476_7351# VPWR 0.156212f
C1906 VPWR _060_ 2.88066f
C1907 VPWR a_9777_2767# 0.190521f
C1908 _080_ VPWR 3.50116f
C1909 net2 _083_ 0.621746f
C1910 counter\[7\] counter\[5\] 0.123194f
C1911 _057_ net7 0.1907f
C1912 _018_ net11 1.60156f
C1913 a_3965_8751# VPWR 0.275213f
C1914 clknet_1_0__leaf_clk _026_ 0.640363f
C1915 _024_ _039_ 0.123357f
C1916 a_2401_8751# a_2842_8863# 0.111047f
C1917 _020_ _033_ 0.522289f
C1918 a_3867_9813# VPWR 0.420123f
C1919 ones[1] _053_ 0.137058f
C1920 _024_ a_5496_9269# 0.231249f
C1921 a_4153_7663# _000_ 0.114647f
C1922 counter\[1\] _055_ 0.226844f
C1923 ones[1] ones[3] 0.371375f
C1924 net2 a_2971_4399# 0.24706f
C1925 _079_ _020_ 0.64168f
C1926 _053_ _055_ 0.242657f
C1927 a_4135_4373# counter\[0\] 0.163031f
C1928 _039_ _086_ 0.185314f
C1929 _049_ net1 0.102595f
C1930 _081_ VPWR 0.336692f
C1931 a_7625_5461# counter\[4\] 0.111904f
C1932 _080_ _023_ 0.187209f
C1933 a_3965_7125# VPWR 0.27379f
C1934 _032_ _027_ 0.291053f
C1935 a_8767_10749# _061_ 0.130378f
C1936 _071_ a_6835_5853# 0.145716f
C1937 _032_ _078_ 0.108688f
C1938 _070_ VPWR 0.29514f
C1939 _038_ _085_ 0.277215f
C1940 a_2295_5461# _010_ 0.101481f
C1941 a_9558_6687# VPWR 0.183627f
C1942 net8 a_4589_3829# 0.169873f
C1943 a_5547_8751# a_5713_8751# 0.966391f
C1944 _014_ _073_ 0.329352f
C1945 _053_ net14 0.290447f
C1946 counter\[1\] _051_ 0.162681f
C1947 _040_ net11 0.200019f
C1948 _030_ clknet_1_1__leaf_clk 0.4999f
C1949 _022_ VPWR 1.67783f
C1950 _053_ _051_ 1.1758f
C1951 a_3394_4917# VPWR 0.192315f
C1952 _016_ VPWR 0.477966f
C1953 _037_ VPWR 0.475818f
C1954 VPWR a_8374_7241# 0.296927f
C1955 _075_ counter\[8\] 0.130767f
C1956 _083_ _073_ 0.29092f
C1957 a_7625_5461# VPWR 0.19847f
C1958 a_7939_9301# a_8105_9301# 0.961627f
C1959 a_9122_2223# counter\[2\] 0.166205f
C1960 net13 net11 1.15219f
C1961 _069_ a_6612_3829# 0.162865f
C1962 a_4526_9813# a_4455_9839# 0.239923f
C1963 _070_ _006_ 0.117927f
C1964 _071_ net1 0.365308f
C1965 counter\[9\] clknet_1_0__leaf_clk 0.264623f
C1966 net7 _061_ 0.227062f
C1967 a_2302_5761# VPWR 0.288521f
C1968 a_4403_6549# a_4694_6849# 0.189515f
C1969 _059_ counter\[1\] 0.364842f
C1970 _048_ _067_ 1.02993f
C1971 net3 _061_ 0.190127f
C1972 a_7987_7828# VPWR 0.254857f
C1973 _039_ _074_ 0.130252f
C1974 _036_ net1 0.287791f
C1975 a_3799_8751# clknet_1_0__leaf_clk 0.299946f
C1976 a_7102_6575# clknet_1_1__leaf_clk 1.74705f
C1977 clk _075_ 0.205306f
C1978 a_6154_8863# VPWR 0.178336f
C1979 net2 a_2787_4949# 0.372244f
C1980 counter\[1\] clknet_1_1__leaf_clk 0.581085f
C1981 _079_ _049_ 0.175275f
C1982 clknet_1_0__leaf_clk _003_ 0.246754f
C1983 _066_ counter\[1\] 1.10194f
C1984 counter\[4\] counter\[6\] 0.278712f
C1985 _009_ _033_ 0.105162f
C1986 net2 net14 2.38473f
C1987 a_4798_5737# VPWR 0.132002f
C1988 _056_ _054_ 0.307119f
C1989 _066_ _053_ 0.176449f
C1990 a_8381_6037# net4 0.368315f
C1991 ones[6] counter\[6\] 0.195496f
C1992 _052_ a_7343_7351# 0.234434f
C1993 rst VGND 0.757091f
C1994 pulse VGND 0.529423f
C1995 ones[2] VGND 0.531794f
C1996 ready VGND 0.5818f
C1997 ones[7] VGND 0.377303f
C1998 ones[6] VGND 0.509771f
C1999 clk VGND 2.67881f
C2000 ones[1] VGND 0.534239f
C2001 ones[5] VGND 0.536071f
C2002 ones[8] VGND 0.57992f
C2003 ones[3] VGND 0.611147f
C2004 ones[0] VGND 0.567651f
C2005 ones[4] VGND 0.436813f
C2006 ones[10] VGND 0.559123f
C2007 ones[9] VGND 0.821373f
C2008 VPWR VGND 0.327472p
C2009 _059_ VGND 2.87205f
C2010 a_10199_2197# VGND 0.384133f
C2011 a_9122_2223# VGND 0.316498f
C2012 a_2511_2223# VGND 0.301339f
C2013 a_1465_2473# VGND 0.378707f
C2014 a_2573_3087# VGND 0.207518f
C2015 a_9648_2741# VGND 0.400385f
C2016 a_8268_2741# VGND 0.34087f
C2017 a_7531_2741# VGND 0.289214f
C2018 a_6375_2767# VGND 0.280197f
C2019 _060_ VGND 0.481499f
C2020 a_4225_2767# VGND 0.370773f
C2021 a_2419_2767# VGND 0.312959f
C2022 _045_ VGND 2.17631f
C2023 a_1761_2999# VGND 0.217798f
C2024 a_4120_3291# VGND 0.226442f
C2025 _032_ VGND 2.02769f
C2026 a_10199_3285# VGND 0.381541f
C2027 a_9011_3285# VGND 0.42363f
C2028 a_8075_3285# VGND 0.30035f
C2029 a_7711_3463# VGND 0.218976f
C2030 a_5731_3311# VGND 0.276649f
C2031 a_3847_3463# VGND 0.253079f
C2032 a_8355_4074# VGND 0.26655f
C2033 a_6612_3829# VGND 0.381857f
C2034 a_4589_3829# VGND 0.290245f
C2035 a_3521_3971# VGND 0.254828f
C2036 a_3421_3855# VGND 0.213288f
C2037 a_10239_4399# VGND 0.223553f
C2038 a_9963_4399# VGND 0.248145f
C2039 a_7607_4765# VGND 0.287772f
C2040 a_7775_4667# VGND 0.350994f
C2041 a_7182_4765# VGND 0.197758f
C2042 a_7350_4511# VGND 0.250219f
C2043 a_6909_4399# VGND 0.328837f
C2044 a_6743_4399# VGND 0.488794f
C2045 a_6135_4765# VGND 0.287573f
C2046 a_6303_4667# VGND 0.357403f
C2047 a_5710_4765# VGND 0.213734f
C2048 a_5878_4511# VGND 0.246324f
C2049 a_5437_4399# VGND 0.30635f
C2050 a_5271_4399# VGND 0.478308f
C2051 _048_ VGND 0.890565f
C2052 a_1407_4399# VGND 0.19535f
C2053 a_5043_4564# VGND 0.219082f
C2054 a_4135_4373# VGND 0.344329f
C2055 a_3137_4765# VGND 0.203576f
C2056 a_2971_4399# VGND 0.250297f
C2057 a_2509_4663# VGND 0.237391f
C2058 a_2409_4445# VGND 0.203485f
C2059 a_1775_4399# VGND 0.224456f
C2060 a_9963_5263# VGND 0.126496f
C2061 a_10136_4943# VGND 0.257984f
C2062 a_9687_4943# VGND 0.255889f
C2063 a_8527_4943# VGND 0.261914f
C2064 a_8695_4917# VGND 0.359157f
C2065 a_8102_4943# VGND 0.206991f
C2066 a_8270_4917# VGND 0.241849f
C2067 a_7829_4949# VGND 0.314173f
C2068 _002_ VGND 0.719866f
C2069 a_7663_4949# VGND 0.509586f
C2070 a_5307_4943# VGND 0.276653f
C2071 a_5475_4917# VGND 0.375795f
C2072 a_4882_4943# VGND 0.209189f
C2073 a_5050_4917# VGND 0.256158f
C2074 a_4609_4949# VGND 0.430776f
C2075 a_4443_4949# VGND 0.48641f
C2076 a_3651_4943# VGND 0.254468f
C2077 a_3819_4917# VGND 0.423249f
C2078 a_3226_4943# VGND 0.200667f
C2079 a_3394_4917# VGND 0.23705f
C2080 a_2953_4949# VGND 0.315546f
C2081 a_2787_4949# VGND 0.488723f
C2082 a_2409_5263# VGND 0.25135f
C2083 _066_ VGND 3.01604f
C2084 _011_ VGND 0.685892f
C2085 a_9735_5639# VGND 0.482557f
C2086 a_9043_5487# VGND 0.256049f
C2087 a_8123_5487# VGND 0.274127f
C2088 a_7625_5461# VGND 0.30768f
C2089 a_6835_5853# VGND 0.251089f
C2090 a_6511_5461# VGND 0.21663f
C2091 a_6335_5461# VGND 0.213869f
C2092 _082_ VGND 1.09613f
C2093 a_5018_5461# VGND 0.353925f
C2094 a_2431_5487# VGND 0.267284f
C2095 a_2502_5461# VGND 0.223586f
C2096 a_2295_5461# VGND 0.521432f
C2097 a_2302_5761# VGND 0.35245f
C2098 a_2011_5461# VGND 0.295367f
C2099 a_1915_5639# VGND 0.395399f
C2100 _081_ VGND 0.286774f
C2101 _037_ VGND 0.700547f
C2102 _057_ VGND 1.20814f
C2103 a_2941_6351# VGND 0.194603f
C2104 _028_ VGND 1.34037f
C2105 a_9739_6005# VGND 0.253671f
C2106 a_9079_6031# VGND 0.27281f
C2107 a_9247_6005# VGND 0.35202f
C2108 a_8654_6031# VGND 0.198649f
C2109 a_8822_6005# VGND 0.244656f
C2110 a_8381_6037# VGND 0.299651f
C2111 _021_ VGND 0.984326f
C2112 a_8215_6037# VGND 0.474557f
C2113 a_7515_6031# VGND 0.274288f
C2114 a_7683_6005# VGND 0.447123f
C2115 a_7090_6031# VGND 0.198034f
C2116 a_7258_6005# VGND 0.241849f
C2117 a_6817_6037# VGND 0.299191f
C2118 a_6651_6037# VGND 0.48674f
C2119 _080_ VGND 0.780011f
C2120 a_4981_6263# VGND 0.215164f
C2121 a_4491_6263# VGND 0.233784f
C2122 a_3851_6005# VGND 0.263489f
C2123 a_2787_6031# VGND 0.340425f
C2124 _046_ VGND 0.404298f
C2125 _043_ VGND 1.26251f
C2126 _047_ VGND 1.17529f
C2127 a_9815_6941# VGND 0.253007f
C2128 a_9983_6843# VGND 0.437665f
C2129 a_9390_6941# VGND 0.197326f
C2130 a_9558_6687# VGND 0.241145f
C2131 a_9117_6575# VGND 0.311595f
C2132 a_8951_6575# VGND 0.487527f
C2133 a_7102_6575# VGND 2.00417f
C2134 _036_ VGND 3.04501f
C2135 a_6060_6549# VGND 0.369048f
C2136 a_2924_6575# VGND 0.227089f
C2137 _065_ VGND 0.957142f
C2138 _006_ VGND 1.15271f
C2139 _018_ VGND 0.44344f
C2140 a_4823_6575# VGND 0.237131f
C2141 a_4894_6549# VGND 0.197031f
C2142 a_4687_6549# VGND 0.498311f
C2143 a_4694_6849# VGND 0.299816f
C2144 a_4403_6549# VGND 0.256696f
C2145 a_4307_6727# VGND 0.33094f
C2146 a_3847_6727# VGND 0.239112f
C2147 _070_ VGND 1.52559f
C2148 a_2734_6575# VGND 0.291723f
C2149 _035_ VGND 2.404f
C2150 a_9661_7439# VGND 0.178561f
C2151 a_9411_7439# VGND 0.103165f
C2152 net2 VGND 1.79914f
C2153 _050_ VGND 1.64399f
C2154 _051_ VGND 1.85527f
C2155 a_8503_7497# VGND 0.256173f
C2156 a_8574_7396# VGND 0.19966f
C2157 a_8374_7241# VGND 0.301798f
C2158 a_8367_7337# VGND 0.480167f
C2159 a_8083_7351# VGND 0.254709f
C2160 a_7987_7351# VGND 0.332294f
C2161 a_7616_7351# VGND 0.220143f
C2162 _005_ VGND 0.471851f
C2163 a_7343_7351# VGND 0.252256f
C2164 a_5823_7119# VGND 0.219681f
C2165 _067_ VGND 0.619425f
C2166 a_4663_7119# VGND 0.253145f
C2167 a_4831_7093# VGND 0.334506f
C2168 a_4238_7119# VGND 0.19384f
C2169 a_4406_7093# VGND 0.236424f
C2170 a_3965_7125# VGND 0.291656f
C2171 _015_ VGND 0.382992f
C2172 a_3799_7125# VGND 0.482155f
C2173 a_3476_7351# VGND 0.198677f
C2174 counter\[10\] VGND 1.13213f
C2175 _049_ VGND 1.39892f
C2176 _014_ VGND 0.493195f
C2177 a_2603_7439# VGND 0.128433f
C2178 _074_ VGND 0.851583f
C2179 a_3203_7351# VGND 0.225982f
C2180 a_2776_7119# VGND 0.246319f
C2181 a_2143_7232# VGND 0.259448f
C2182 _085_ VGND 1.7836f
C2183 a_9815_8029# VGND 0.254513f
C2184 a_9983_7931# VGND 0.35449f
C2185 a_9390_8029# VGND 0.194813f
C2186 a_9558_7775# VGND 0.24121f
C2187 a_9117_7663# VGND 0.311364f
C2188 _020_ VGND 1.1992f
C2189 a_8951_7663# VGND 0.495776f
C2190 a_7987_7828# VGND 0.245758f
C2191 net6 VGND 1.9055f
C2192 a_7263_7637# VGND 0.348365f
C2193 a_5433_7637# VGND 1.98941f
C2194 a_4663_8029# VGND 0.257066f
C2195 a_4831_7931# VGND 0.418554f
C2196 a_4238_8029# VGND 0.193124f
C2197 a_4406_7775# VGND 0.239857f
C2198 a_3965_7663# VGND 0.327118f
C2199 a_3799_7663# VGND 0.486591f
C2200 a_3099_8029# VGND 0.270192f
C2201 a_3267_7931# VGND 0.369971f
C2202 a_2674_8029# VGND 0.233091f
C2203 a_2842_7775# VGND 0.264665f
C2204 a_2401_7663# VGND 0.347038f
C2205 a_2235_7663# VGND 0.522854f
C2206 a_2007_7828# VGND 0.249001f
C2207 a_8863_8527# VGND 0.219746f
C2208 _010_ VGND 0.78645f
C2209 _056_ VGND 2.30234f
C2210 _073_ VGND 0.830201f
C2211 _000_ VGND 0.654088f
C2212 net1 VGND 2.32668f
C2213 a_9926_8181# VGND 0.307779f
C2214 a_9503_8207# VGND 0.218827f
C2215 _079_ VGND 1.18052f
C2216 _078_ VGND 2.33271f
C2217 a_8727_8181# VGND 0.262242f
C2218 a_7239_8207# VGND 0.266465f
C2219 a_7407_8181# VGND 0.451366f
C2220 a_6814_8207# VGND 0.202421f
C2221 a_6982_8181# VGND 0.243744f
C2222 a_6541_8213# VGND 0.298505f
C2223 _008_ VGND 0.636644f
C2224 a_6375_8213# VGND 0.483152f
C2225 clknet_0_clk VGND 2.33677f
C2226 a_3593_8181# VGND 2.00425f
C2227 a_2879_8207# VGND 0.273773f
C2228 _054_ VGND 0.695229f
C2229 _044_ VGND 2.81787f
C2230 _055_ VGND 0.905885f
C2231 a_10239_8751# VGND 0.265955f
C2232 a_9687_8751# VGND 0.217446f
C2233 a_9411_8751# VGND 0.230621f
C2234 a_7833_8903# VGND 0.242522f
C2235 a_6411_9117# VGND 0.292429f
C2236 a_6579_9019# VGND 0.507146f
C2237 a_5986_9117# VGND 0.213825f
C2238 a_6154_8863# VGND 0.259721f
C2239 a_5713_8751# VGND 0.328376f
C2240 _001_ VGND 2.7776f
C2241 a_5547_8751# VGND 0.466213f
C2242 _016_ VGND 0.612904f
C2243 a_5271_8751# VGND 0.211924f
C2244 _033_ VGND 0.632748f
C2245 a_4663_9117# VGND 0.259359f
C2246 a_4831_9019# VGND 0.336642f
C2247 a_4238_9117# VGND 0.206382f
C2248 a_4406_8863# VGND 0.250252f
C2249 a_3965_8751# VGND 0.304513f
C2250 _012_ VGND 1.78482f
C2251 a_3799_8751# VGND 0.500842f
C2252 a_3099_9117# VGND 0.277358f
C2253 a_3267_9019# VGND 0.358619f
C2254 a_2674_9117# VGND 0.244222f
C2255 a_2842_8863# VGND 0.276746f
C2256 a_2401_8751# VGND 0.345774f
C2257 a_2235_8751# VGND 0.548822f
C2258 _013_ VGND 0.541218f
C2259 net14 VGND 2.4358f
C2260 _042_ VGND 1.48931f
C2261 _026_ VGND 0.452907f
C2262 counter\[9\] VGND 3.97321f
C2263 a_10103_9514# VGND 0.240812f
C2264 a_9551_9527# VGND 0.245874f
C2265 a_8803_9295# VGND 0.276703f
C2266 a_8971_9269# VGND 0.356027f
C2267 a_8378_9295# VGND 0.209164f
C2268 a_8546_9269# VGND 0.255851f
C2269 a_8105_9301# VGND 0.324271f
C2270 _022_ VGND 0.743005f
C2271 a_7939_9301# VGND 0.513495f
C2272 clknet_1_1__leaf_clk VGND 3.95119f
C2273 _040_ VGND 0.833938f
C2274 _041_ VGND 0.437873f
C2275 a_5871_9527# VGND 0.267044f
C2276 a_5496_9269# VGND 0.253205f
C2277 net7 VGND 2.18383f
C2278 _009_ VGND 0.319397f
C2279 a_4363_9673# VGND 0.242551f
C2280 a_4434_9572# VGND 0.196486f
C2281 a_4234_9417# VGND 0.298321f
C2282 a_4227_9513# VGND 0.489386f
C2283 a_3943_9527# VGND 0.258424f
C2284 a_3847_9527# VGND 0.352774f
C2285 _052_ VGND 1.60879f
C2286 a_3300_9269# VGND 0.332492f
C2287 _053_ VGND 4.70496f
C2288 _076_ VGND 2.64432f
C2289 _075_ VGND 4.00525f
C2290 _077_ VGND 0.559357f
C2291 _004_ VGND 1.28767f
C2292 _062_ VGND 0.517851f
C2293 a_10103_9991# VGND 0.257423f
C2294 a_9779_9839# VGND 0.241842f
C2295 _064_ VGND 1.58568f
C2296 a_6324_10029# VGND 0.288755f
C2297 a_5513_10089# VGND 0.329389f
C2298 counter\[3\] VGND 2.16401f
C2299 _003_ VGND 0.635499f
C2300 net12 VGND 6.54231f
C2301 a_4455_9839# VGND 0.240169f
C2302 a_4526_9813# VGND 0.197548f
C2303 a_4319_9813# VGND 0.4851f
C2304 a_4326_10113# VGND 0.299908f
C2305 a_4035_9813# VGND 0.276335f
C2306 a_3867_9813# VGND 0.459816f
C2307 _063_ VGND 0.655318f
C2308 a_3479_10004# VGND 0.262927f
C2309 a_2271_10205# VGND 0.300695f
C2310 a_2439_10107# VGND 0.537251f
C2311 a_1846_10205# VGND 0.221206f
C2312 a_2014_9951# VGND 0.265308f
C2313 a_1573_9839# VGND 0.454954f
C2314 _019_ VGND 0.647811f
C2315 a_1407_9839# VGND 0.560011f
C2316 clknet_1_0__leaf_clk VGND 4.64197f
C2317 _068_ VGND 1.58845f
C2318 net9 VGND 6.88615f
C2319 _034_ VGND 0.914748f
C2320 _058_ VGND 1.4918f
C2321 _084_ VGND 0.863911f
C2322 a_10239_10383# VGND 0.219801f
C2323 net8 VGND 4.02803f
C2324 a_9963_10383# VGND 0.244545f
C2325 net4 VGND 1.26275f
C2326 a_8767_10749# VGND 0.296047f
C2327 _061_ VGND 5.92109f
C2328 counter\[6\] VGND 2.24659f
C2329 counter\[4\] VGND 2.36668f
C2330 counter\[5\] VGND 2.91211f
C2331 a_8091_10615# VGND 0.274625f
C2332 counter\[2\] VGND 1.9989f
C2333 counter\[1\] VGND 5.14823f
C2334 counter\[0\] VGND 5.37383f
C2335 _083_ VGND 3.4741f
C2336 net3 VGND 6.38788f
C2337 net5 VGND 2.11089f
C2338 a_7729_10927# VGND 0.120944f
C2339 a_7479_10927# VGND 0.241885f
C2340 a_7197_10927# VGND 0.133165f
C2341 _072_ VGND 2.76201f
C2342 _039_ VGND 1.74718f
C2343 _007_ VGND 0.965425f
C2344 _017_ VGND 0.611544f
C2345 _030_ VGND 0.772848f
C2346 a_10134_10927# VGND 0.276684f
C2347 counter\[8\] VGND 2.49678f
C2348 a_9687_10927# VGND 0.244882f
C2349 net13 VGND 1.82078f
C2350 _031_ VGND 3.93171f
C2351 net10 VGND 2.60709f
C2352 net11 VGND 4.6317f
C2353 counter\[7\] VGND 7.89787f
C2354 _069_ VGND 4.4444f
C2355 _071_ VGND 0.774167f
C2356 a_6979_10901# VGND 0.252709f
C2357 _038_ VGND 1.57063f
C2358 a_5503_11092# VGND 0.261944f
C2359 a_4901_11191# VGND 0.240285f
C2360 _029_ VGND 0.801813f
C2361 a_4801_10973# VGND 0.212498f
C2362 _025_ VGND 0.838692f
C2363 _024_ VGND 5.79771f
C2364 _027_ VGND 3.09769f
C2365 a_1773_11191# VGND 0.253112f
C2366 _023_ VGND 3.70689f
C2367 a_1673_10973# VGND 0.214109f
C2368 _086_ VGND 5.49993f
.ends

