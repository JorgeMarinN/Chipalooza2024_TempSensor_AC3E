magic
tech sky130A
timestamp 1713593032
<< error_s >>
rect 5 196 95 830
rect 4 95 196 196
rect 4 86 389 95
rect 4 14 396 86
rect 4 5 389 14
rect 4 4 196 5
use vias_gen$16  vias_gen$16_0
timestamp 1713593032
transform 1 0 0 0 1 0
box 0 0 100 100
use vias_gen$18  vias_gen$18_0
timestamp 1713593032
transform 1 0 0 0 1 0
box 0 0 400 100
use vias_gen$19  vias_gen$19_0
timestamp 1713593032
transform 1 0 0 0 1 0
box 0 0 400 100
use vias_gen$21  vias_gen$21_0
timestamp 1713593032
transform 1 0 0 0 1 0
box 0 0 100 100
use vias_gen$22  vias_gen$22_0
timestamp 1713593032
transform 1 0 0 0 1 0
box 0 0 200 200
use vias_gen$23  vias_gen$23_0
timestamp 1713593032
transform 1 0 0 0 1 0
box -13 -13 113 1013
use vias_gen$24  vias_gen$24_0
timestamp 1713593032
transform 1 0 0 0 1 0
box 0 0 150 200
use vias_gen$25  vias_gen$25_0
timestamp 1713593032
transform 1 0 0 0 1 0
box 0 0 200 200
use vias_gen$26  vias_gen$26_0
timestamp 1713593032
transform 1 0 0 0 1 0
box 0 0 100 200
<< end >>
