magic
tech sky130A
magscale 1 2
timestamp 1713591521
<< pwell >>
rect -729 1286 729 1372
rect -729 -1372 729 -1286
<< psubdiff >>
rect -703 1312 -595 1346
rect -561 1312 -527 1346
rect -493 1312 -459 1346
rect -425 1312 -391 1346
rect -357 1312 -323 1346
rect -289 1312 -255 1346
rect -221 1312 -187 1346
rect -153 1312 -119 1346
rect -85 1312 -51 1346
rect -17 1312 17 1346
rect 51 1312 85 1346
rect 119 1312 153 1346
rect 187 1312 221 1346
rect 255 1312 289 1346
rect 323 1312 357 1346
rect 391 1312 425 1346
rect 459 1312 493 1346
rect 527 1312 561 1346
rect 595 1312 703 1346
rect -703 -1346 -595 -1312
rect -561 -1346 -527 -1312
rect -493 -1346 -459 -1312
rect -425 -1346 -391 -1312
rect -357 -1346 -323 -1312
rect -289 -1346 -255 -1312
rect -221 -1346 -187 -1312
rect -153 -1346 -119 -1312
rect -85 -1346 -51 -1312
rect -17 -1346 17 -1312
rect 51 -1346 85 -1312
rect 119 -1346 153 -1312
rect 187 -1346 221 -1312
rect 255 -1346 289 -1312
rect 323 -1346 357 -1312
rect 391 -1346 425 -1312
rect 459 -1346 493 -1312
rect 527 -1346 561 -1312
rect 595 -1346 703 -1312
<< psubdiffcont >>
rect -595 1312 -561 1346
rect -527 1312 -493 1346
rect -459 1312 -425 1346
rect -391 1312 -357 1346
rect -323 1312 -289 1346
rect -255 1312 -221 1346
rect -187 1312 -153 1346
rect -119 1312 -85 1346
rect -51 1312 -17 1346
rect 17 1312 51 1346
rect 85 1312 119 1346
rect 153 1312 187 1346
rect 221 1312 255 1346
rect 289 1312 323 1346
rect 357 1312 391 1346
rect 425 1312 459 1346
rect 493 1312 527 1346
rect 561 1312 595 1346
rect -595 -1346 -561 -1312
rect -527 -1346 -493 -1312
rect -459 -1346 -425 -1312
rect -391 -1346 -357 -1312
rect -323 -1346 -289 -1312
rect -255 -1346 -221 -1312
rect -187 -1346 -153 -1312
rect -119 -1346 -85 -1312
rect -51 -1346 -17 -1312
rect 17 -1346 51 -1312
rect 85 -1346 119 -1312
rect 153 -1346 187 -1312
rect 221 -1346 255 -1312
rect 289 -1346 323 -1312
rect 357 -1346 391 -1312
rect 425 -1346 459 -1312
rect 493 -1346 527 -1312
rect 561 -1346 595 -1312
<< xpolycontact >>
rect -573 784 573 1216
rect -573 -1216 573 -784
<< ppolyres >>
rect -573 -784 573 784
<< locali >>
rect -703 1312 -595 1346
rect -561 1312 -527 1346
rect -493 1312 -459 1346
rect -425 1312 -391 1346
rect -357 1312 -323 1346
rect -289 1312 -255 1346
rect -221 1312 -187 1346
rect -153 1312 -119 1346
rect -85 1312 -51 1346
rect -17 1312 17 1346
rect 51 1312 85 1346
rect 119 1312 153 1346
rect 187 1312 221 1346
rect 255 1312 289 1346
rect 323 1312 357 1346
rect 391 1312 425 1346
rect 459 1312 493 1346
rect 527 1312 561 1346
rect 595 1312 703 1346
rect -703 -1346 -595 -1312
rect -561 -1346 -527 -1312
rect -493 -1346 -459 -1312
rect -425 -1346 -391 -1312
rect -357 -1346 -323 -1312
rect -289 -1346 -255 -1312
rect -221 -1346 -187 -1312
rect -153 -1346 -119 -1312
rect -85 -1346 -51 -1312
rect -17 -1346 17 -1312
rect 51 -1346 85 -1312
rect 119 -1346 153 -1312
rect 187 -1346 221 -1312
rect 255 -1346 289 -1312
rect 323 -1346 357 -1312
rect 391 -1346 425 -1312
rect 459 -1346 493 -1312
rect 527 -1346 561 -1312
rect 595 -1346 703 -1312
<< viali >>
rect -557 802 557 1196
rect -557 -1197 557 -803
<< metal1 >>
rect -569 1196 569 1204
rect -569 802 -557 1196
rect 557 802 569 1196
rect -569 795 569 802
rect -569 -803 569 -795
rect -569 -1197 -557 -803
rect 557 -1197 569 -803
rect -569 -1204 569 -1197
<< properties >>
string FIXED_BBOX -686 -1329 686 1329
<< end >>
