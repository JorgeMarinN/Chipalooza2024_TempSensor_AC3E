magic
tech sky130A
magscale 1 2
timestamp 1713593032
<< pwell >>
rect -26 -26 226 226
<< psubdiff >>
rect 0 151 200 200
rect 0 49 49 151
rect 151 49 200 151
rect 0 0 200 49
<< psubdiffcont >>
rect 49 49 151 151
<< locali >>
rect 0 153 200 200
rect 0 47 47 153
rect 153 47 200 153
rect 0 0 200 47
<< viali >>
rect 47 151 153 153
rect 47 49 49 151
rect 49 49 151 151
rect 151 49 153 151
rect 47 47 153 49
<< metal1 >>
rect 0 190 200 200
rect 0 10 10 190
rect 190 10 200 190
rect 0 0 200 10
<< via1 >>
rect 10 153 190 190
rect 10 47 47 153
rect 47 47 153 153
rect 153 47 190 153
rect 10 10 190 47
<< metal2 >>
rect 0 190 200 200
rect 0 10 10 190
rect 190 10 200 190
rect 0 0 200 10
<< via2 >>
rect 32 32 168 168
<< metal3 >>
rect 0 168 200 200
rect 0 32 32 168
rect 168 32 200 168
rect 0 0 200 32
<< end >>
