magic
tech sky130A
timestamp 1713593032
<< metal4 >>
rect -40 959 1322 1040
rect -40 841 1181 959
rect 1299 841 1322 959
rect -40 799 1322 841
rect -40 681 1181 799
rect 1299 681 1322 799
rect -40 639 1322 681
rect -40 521 1181 639
rect 1299 521 1322 639
rect -40 479 1322 521
rect -40 361 1181 479
rect 1299 361 1322 479
rect -40 319 1322 361
rect -40 201 1181 319
rect 1299 201 1322 319
rect -40 159 1322 201
rect -40 41 1181 159
rect 1299 41 1322 159
rect -40 -40 1322 41
<< via4 >>
rect 1181 841 1299 959
rect 1181 681 1299 799
rect 1181 521 1299 639
rect 1181 361 1299 479
rect 1181 201 1299 319
rect 1181 41 1299 159
<< mimcap2 >>
rect 0 959 1000 1000
rect 0 41 41 959
rect 959 41 1000 959
rect 0 0 1000 41
<< mimcap2contact >>
rect 41 41 959 959
<< metal5 >>
rect 8 959 992 992
rect 8 41 41 959
rect 959 41 992 959
rect 8 8 992 41
rect 1160 959 1320 1034
rect 1160 841 1181 959
rect 1299 841 1320 959
rect 1160 799 1320 841
rect 1160 681 1181 799
rect 1299 681 1320 799
rect 1160 639 1320 681
rect 1160 521 1181 639
rect 1299 521 1320 639
rect 1160 479 1320 521
rect 1160 361 1181 479
rect 1299 361 1320 479
rect 1160 319 1320 361
rect 1160 201 1181 319
rect 1299 201 1320 319
rect 1160 159 1320 201
rect 1160 41 1181 159
rect 1299 41 1320 159
rect 1160 -34 1320 41
<< end >>
