* NGSPICE file created from SDC_pex.ext - technology: sky130A

.subckt SDC_pex VDD VSS N2_R DOUT
X0 N3_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 N3_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y INTERNAL_SDC_0.N2_S VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6 VSS VSS VSS sky130_fd_pr__res_high_po_5p73 l=8
X7 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 SENS_IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X8 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X11 VSS a_n10739_n4824# a_n10642_n4576# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X12 INTERNAL_SDC_0.OSC_PGATE_1.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X13 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X14 VDD SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X15 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X16 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X18 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VDD SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X20 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 SENS_IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X23 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y N2_R VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_n10312_n3776# a_n10739_n4824# DOUT VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X25 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 REF_IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 N3_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X27 VDD SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X28 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X29 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X31 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X32 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X35 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X36 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X37 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X38 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 VSS REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X40 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X41 INTERNAL_SDC_0.OSC_PGATE_0.VIN VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X42 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X43 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X44 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X45 SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y INTERNAL_SDC_0.OSC_PGATE_0.VIN VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X46 VDD INTERNAL_SDC_0.N2_S a_n10642_n3576# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X47 INTERNAL_SDC_0.OSC_PGATE_1.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y VDD VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X48 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X49 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X50 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X51 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 REF_IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X52 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X53 INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y DOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X54 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X55 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X56 VDD REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X57 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X58 INTERNAL_SDC_0.OSC_PGATE_0.VIN DOUT SENS_IN VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X59 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 REF_IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X60 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X61 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X62 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X63 SENS_IN VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X64 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X65 INTERNAL_SDC_0.OSC_PGATE_1.VIN INTERNAL_SDC_0.OSC_PGATE_1.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y REF_IN VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X66 VDD SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X67 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X68 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X69 INTERNAL_SDC_0.OSC_PGATE_0.VIN INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y SENS_IN VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X70 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X71 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X72 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X73 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X74 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X75 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 REF_IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X76 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X77 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X78 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X79 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X80 VSS SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X81 REF_IN INTERNAL_SDC_0.OSC_PGATE_1.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y INTERNAL_SDC_0.OSC_PGATE_1.VIN VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X82 SENS_IN VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X83 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X84 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X85 N3_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X86 N3_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X87 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X88 N3_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X89 N2_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X90 VDD VDD VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X91 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X92 INTERNAL_SDC_0.DFF_0.ND a_n10642_n4576# a_n10312_n4576# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X93 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X94 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y N2_R VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X95 INTERNAL_SDC_0.OSC_PGATE_1.VIN INTERNAL_SDC_0.OSC_PGATE_1.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y REF_IN VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X96 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X97 N3_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X98 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X99 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X100 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X101 N3_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X102 a_n10739_n4824# INTERNAL_SDC_0.N2_S VSS VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X103 DOUT INTERNAL_SDC_0.DFF_0.ND VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X104 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X105 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X106 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X107 VSS VSS VSS sky130_fd_pr__res_high_po_5p73 l=8
X108 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X109 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X110 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X111 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X112 INTERNAL_SDC_0.OSC_PGATE_0.VIN INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y SENS_IN VDD sky130_fd_pr__pfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X113 INTERNAL_SDC_0.OSC_PGATE_1.VIN VDD REF_IN VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X114 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X115 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X116 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X117 VSS SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X118 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X119 VDD VDD VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X120 VSS SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X121 INTERNAL_SDC_0.N2_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X122 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 REF_IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X123 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X124 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X125 VDD VDD VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X126 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X127 VSS REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X128 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X129 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X130 VSS SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X131 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X132 INTERNAL_SDC_0.OSC_PGATE_1.VIN VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X133 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X134 N3_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X135 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X136 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X137 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X138 N3_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X139 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X140 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X141 REF_IN VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X142 VDD VDD VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X143 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X144 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X145 VDD SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X146 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X147 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 SENS_IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X148 SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y INTERNAL_SDC_0.OSC_PGATE_0.VIN VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X149 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X150 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y INTERNAL_SDC_0.N2_S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X151 VDD REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X152 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X153 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X154 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X155 SENS_IN N3_S VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X156 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X157 VSS REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X158 N3_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X159 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X160 a_n10642_n4576# N2_R a_n10642_n4776# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X161 N2_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X162 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X163 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X164 VSS SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X165 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X166 VDD VDD VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X167 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X168 a_n10642_n3576# N2_R a_n10739_n4824# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X169 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X170 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X171 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X172 N3_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X173 VDD VDD VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X174 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X175 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X176 DOUT INTERNAL_SDC_0.DFF_0.ND VSS VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X177 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X178 REF_IN VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X179 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X180 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X181 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X182 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 SENS_IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X183 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X184 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X185 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X186 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X187 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X188 SENS_IN N3_S VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X189 N3_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X190 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X191 N3_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X192 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X193 SENS_IN N3_S VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X194 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X195 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X196 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X197 INTERNAL_SDC_0.OSC_PGATE_1.VIN VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X198 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X199 N3_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X200 REF_IN N3_R VSS sky130_fd_pr__res_high_po_5p73 l=8
X201 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X202 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X203 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X204 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X205 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X206 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X207 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X208 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X209 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X210 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X211 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X212 N3_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X213 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X214 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X215 VSS REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X216 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X217 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 REF_IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X218 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X219 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 SENS_IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X220 INTERNAL_SDC_0.OSC_PGATE_0.VIN INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y SENS_IN VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X221 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X222 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X223 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 SENS_IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X224 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X225 a_n10312_n4576# N2_R VSS VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X226 VSS REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X227 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X228 REF_IN VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X229 INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y DOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X230 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X231 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X232 N3_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X233 REF_IN INTERNAL_SDC_0.OSC_PGATE_1.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y INTERNAL_SDC_0.OSC_PGATE_1.VIN VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X234 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X235 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X236 N3_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X237 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 REF_IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X238 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X239 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X240 SENS_IN DOUT INTERNAL_SDC_0.OSC_PGATE_0.VIN VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X241 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X242 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X243 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X244 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X245 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X246 VSS N2_R a_n10312_n3776# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X247 VDD DOUT INTERNAL_SDC_0.DFF_0.ND VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X248 VDD REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X249 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X250 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X251 N3_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X252 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 SENS_IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X253 VSS SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X254 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X255 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X256 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X257 SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y INTERNAL_SDC_0.OSC_PGATE_0.VIN VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X258 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X259 SENS_IN N3_S VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X260 SENS_IN N3_S VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X261 INTERNAL_SDC_0.OSC_PGATE_1.VIN INTERNAL_SDC_0.OSC_PGATE_1.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y REF_IN VDD sky130_fd_pr__pfet_01v8 ad=0.31 pd=2.62 as=0.165 ps=1.33 w=1 l=0.15
X262 SENS_IN N3_S VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X263 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X264 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X265 SENS_IN N3_S VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X266 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 SENS_IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X267 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X268 INTERNAL_SDC_0.N2_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X269 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 REF_IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X270 N3_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X271 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X272 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 SENS_IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X273 N3_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X274 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X275 VDD REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X276 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X277 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X278 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X279 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X280 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X281 REF_IN INTERNAL_SDC_0.OSC_PGATE_1.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y INTERNAL_SDC_0.OSC_PGATE_1.VIN VDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X282 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X283 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X284 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X285 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X286 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X287 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X288 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X289 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X290 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 REF_IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X291 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X292 SENS_IN N3_S VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X293 SENS_IN N3_S VDD sky130_fd_pr__res_iso_pw w=20 l=30.5
X294 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X295 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 SENS_IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X296 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X297 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X298 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X299 VSS REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X300 N3_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X301 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X302 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X303 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X304 a_n10642_n4776# a_n10739_n4824# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X305 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 REF_IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X306 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X307 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X308 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X309 VSS DOUT INTERNAL_SDC_0.DFF_0.ND VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X310 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X311 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X312 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 REF_IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X313 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X314 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__cap_mim_m3_2 l=10 w=10
X315 INTERNAL_SDC_0.OSC_PGATE_0.VIN VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X316 N3_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X317 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X318 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X319 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X320 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X321 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X322 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X323 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X324 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X325 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X326 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X327 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X328 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X329 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 SENS_IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X330 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X331 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X332 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X333 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 SENS_IN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X334 VDD SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X335 VDD REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X336 REF_IN VDD INTERNAL_SDC_0.OSC_PGATE_1.VIN VSS sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.31 ps=2.62 w=1 l=0.15
X337 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X338 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 REF_IN VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X339 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X340 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X341 SENS_IN VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X342 N3_R INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X343 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X344 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X345 VSS INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X346 VDD REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X347 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X348 VDD INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X349 VSS INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X350 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X351 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X352 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X353 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
C0 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out 0.908329f
C1 INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y SENS_IN 0.243798f
C2 REF_IN INTERNAL_SDC_0.OSC_PGATE_1.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y 0.245165f
C3 SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out 0.74966f
C4 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out 0.906047f
C5 a_n10642_n4776# a_n10642_n4576# 0.252453f
C6 REF_IN VDD 1.67939f
C7 REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out 0.74966f
C8 REF_IN INTERNAL_SDC_0.OSC_PGATE_1.VIN 1.87951f
C9 INTERNAL_SDC_0.N2_S N3_S 0.386303f
C10 INTERNAL_SDC_0.DFF_0.ND a_n10642_n4576# 0.157962f
C11 a_n10312_n4576# a_n10642_n4576# 0.17245f
C12 N3_R N2_R 0.370157f
C13 DOUT INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y 0.129257f
C14 N3_R VDD 2.13277f
C15 SENS_IN N3_S 12.787f
C16 INTERNAL_SDC_0.OSC_PGATE_0.VIN SENS_IN 1.87885f
C17 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VDD 3.92679f
C18 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y 0.354794f
C19 DOUT INTERNAL_SDC_0.DFF_0.ND 0.304507f
C20 a_n10642_n4776# VDD 0.222652f
C21 INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y VDD 1.37268f
C22 SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 1.66372f
C23 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out 3.19892f
C24 INTERNAL_SDC_0.DFF_0.ND a_n10739_n4824# 0.11706f
C25 INTERNAL_SDC_0.DFF_0.ND N2_R 0.158287f
C26 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out 0.906047f
C27 INTERNAL_SDC_0.DFF_0.ND VDD 0.674592f
C28 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y N2_R 0.11977f
C29 REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT 0.74966f
C30 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y VDD 0.354794f
C31 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT N3_S 0.887654f
C32 DOUT INTERNAL_SDC_0.OSC_PGATE_0.VIN 0.15133f
C33 INTERNAL_SDC_0.N2_S VDD 2.18027f
C34 DOUT SENS_IN 0.348221f
C35 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VDD 3.19675f
C36 SENS_IN INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT 0.74966f
C37 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 0.906047f
C38 N3_S VDD 80.8389f
C39 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT N3_R 0.887654f
C40 INTERNAL_SDC_0.OSC_PGATE_0.VIN VDD 0.829031f
C41 SENS_IN VDD 80.5525f
C42 VDD INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 3.19675f
C43 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VDD 3.19892f
C44 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out 0.906047f
C45 a_n10642_n4576# a_n10739_n4824# 0.1448f
C46 REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 1.66372f
C47 a_n10312_n3776# DOUT 0.162484f
C48 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out SENS_IN 0.74966f
C49 a_n10642_n3576# a_n10739_n4824# 0.255061f
C50 N2_R a_n10642_n4576# 0.475838f
C51 a_n10642_n4576# VDD 0.109572f
C52 a_n10642_n3576# VDD 0.223093f
C53 a_n10312_n3776# a_n10739_n4824# 0.213834f
C54 REF_IN SENS_IN 8.17084f
C55 REF_IN INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out 0.74966f
C56 DOUT a_n10739_n4824# 0.289294f
C57 DOUT N2_R 0.194525f
C58 DOUT VDD 1.26612f
C59 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VDD 3.92679f
C60 INTERNAL_SDC_0.N2_S INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y 0.126003f
C61 INTERNAL_SDC_0.OSC_PGATE_1.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y VDD 1.51486f
C62 a_n10312_n4576# INTERNAL_SDC_0.DFF_0.ND 0.162484f
C63 N2_R a_n10739_n4824# 0.530612f
C64 INTERNAL_SDC_0.OSC_PGATE_1.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y INTERNAL_SDC_0.OSC_PGATE_1.VIN 0.261217f
C65 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT 0.908329f
C66 a_n10739_n4824# VDD 0.782611f
C67 N2_R VDD 1.89719f
C68 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VDD 3.19892f
C69 INTERNAL_SDC_0.OSC_PGATE_1.VIN VDD 0.957623f
C70 INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y INTERNAL_SDC_0.OSC_PGATE_0.VIN 0.261021f
C71 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VDD 3.19892f
C72 N2_R VSS 10.2263f
C73 DOUT VSS 4.83678f
C74 VDD VSS 2.10313p
C75 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y VSS 0.462218f
C76 N3_R VSS 6.61484f
C77 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.INVandCAP_0[3].VOUT VSS 65.84f
C78 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x2_out VSS 64.070206f
C79 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.x1_out VSS 64.0533f
C80 INTERNAL_SDC_0.OSC_PGATE_1.OSC_0.N1 VSS 64.0406f
C81 INTERNAL_SDC_0.OSC_PGATE_1.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y VSS 0.622583f
C82 REF_IN VSS 59.757496f
C83 INTERNAL_SDC_0.OSC_PGATE_1.VIN VSS 23.837f
C84 a_n10312_n4576# VSS 0.242922f
C85 a_n10642_n4576# VSS 0.786451f
C86 INTERNAL_SDC_0.DFF_0.ND VSS 0.389686f
C87 a_n10312_n3776# VSS 0.239496f
C88 a_n10739_n4824# VSS 1.21396f
C89 INTERNAL_SDC_0.OSC_PGATE_0.VIN VSS 23.788f
C90 INTERNAL_SDC_0.OSC_PGATE_0.PASSGATE_0.sky130_fd_sc_hd__inv_1$1_0.Y VSS 0.628215f
C91 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x2_out VSS 64.070206f
C92 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.x1_out VSS 64.0533f
C93 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.N1 VSS 64.0406f
C94 INTERNAL_SDC_0.N2_S VSS 8.590549f
C95 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.BUFFMIN_0.sky130_fd_sc_hd__inv_1_0.Y VSS 0.462218f
C96 INTERNAL_SDC_0.OSC_PGATE_0.OSC_0.INVandCAP_0[3].VOUT VSS 65.8343f
C97 N3_S VSS 43.1455f
C98 SENS_IN VSS 94.6087f
.ends

