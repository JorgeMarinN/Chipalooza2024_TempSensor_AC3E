magic
tech sky130A
magscale 1 2
timestamp 1713593032
<< viali >>
rect 1593 11305 1627 11339
rect 4077 11305 4111 11339
rect 8493 11305 8527 11339
rect 3341 11237 3375 11271
rect 5273 11237 5307 11271
rect 8769 11237 8803 11271
rect 2421 11169 2455 11203
rect 2605 11169 2639 11203
rect 2697 11169 2731 11203
rect 2789 11169 2823 11203
rect 1501 11101 1535 11135
rect 2881 11101 2915 11135
rect 4353 11101 4387 11135
rect 4445 11101 4479 11135
rect 5733 11101 5767 11135
rect 5825 11101 5859 11135
rect 8309 11101 8343 11135
rect 8585 11101 8619 11135
rect 8953 11101 8987 11135
rect 3065 11033 3099 11067
rect 4629 11033 4663 11067
rect 5549 11033 5583 11067
rect 9198 11033 9232 11067
rect 3525 10965 3559 10999
rect 4261 10965 4295 10999
rect 10333 10965 10367 10999
rect 1869 10761 1903 10795
rect 7205 10761 7239 10795
rect 7389 10761 7423 10795
rect 8033 10761 8067 10795
rect 8493 10761 8527 10795
rect 2481 10693 2515 10727
rect 2697 10693 2731 10727
rect 9290 10693 9324 10727
rect 1501 10625 1535 10659
rect 1777 10625 1811 10659
rect 2881 10625 2915 10659
rect 3065 10625 3099 10659
rect 7481 10625 7515 10659
rect 7849 10625 7883 10659
rect 8309 10625 8343 10659
rect 8585 10625 8619 10659
rect 8769 10625 8803 10659
rect 9045 10625 9079 10659
rect 1986 10557 2020 10591
rect 7113 10557 7147 10591
rect 7573 10557 7607 10591
rect 2145 10421 2179 10455
rect 2329 10421 2363 10455
rect 2513 10421 2547 10455
rect 2973 10421 3007 10455
rect 7757 10421 7791 10455
rect 8953 10421 8987 10455
rect 10425 10421 10459 10455
rect 4537 10217 4571 10251
rect 4721 10217 4755 10251
rect 9229 10217 9263 10251
rect 3157 10149 3191 10183
rect 2605 10081 2639 10115
rect 3617 10081 3651 10115
rect 8585 10081 8619 10115
rect 1685 10013 1719 10047
rect 2881 10013 2915 10047
rect 3433 10013 3467 10047
rect 3801 10013 3835 10047
rect 4077 10013 4111 10047
rect 4813 10013 4847 10047
rect 4997 10013 5031 10047
rect 6009 10013 6043 10047
rect 6285 10013 6319 10047
rect 6561 10013 6595 10047
rect 4353 9945 4387 9979
rect 6806 9945 6840 9979
rect 9873 9945 9907 9979
rect 9965 9945 9999 9979
rect 10241 9945 10275 9979
rect 1501 9877 1535 9911
rect 2789 9877 2823 9911
rect 2973 9877 3007 9911
rect 3249 9877 3283 9911
rect 3893 9877 3927 9911
rect 4261 9877 4295 9911
rect 4553 9877 4587 9911
rect 4905 9877 4939 9911
rect 6101 9877 6135 9911
rect 6469 9877 6503 9911
rect 7941 9877 7975 9911
rect 9689 9877 9723 9911
rect 10057 9877 10091 9911
rect 2513 9673 2547 9707
rect 6009 9673 6043 9707
rect 3249 9605 3283 9639
rect 4914 9605 4948 9639
rect 8217 9605 8251 9639
rect 8953 9605 8987 9639
rect 1869 9537 1903 9571
rect 2329 9537 2363 9571
rect 6009 9537 6043 9571
rect 6193 9537 6227 9571
rect 7501 9537 7535 9571
rect 9597 9537 9631 9571
rect 9781 9537 9815 9571
rect 9965 9537 9999 9571
rect 10241 9537 10275 9571
rect 5181 9469 5215 9503
rect 7757 9469 7791 9503
rect 2881 9401 2915 9435
rect 3433 9401 3467 9435
rect 8585 9401 8619 9435
rect 8769 9401 8803 9435
rect 9321 9401 9355 9435
rect 9505 9401 9539 9435
rect 2053 9333 2087 9367
rect 3249 9333 3283 9367
rect 3801 9333 3835 9367
rect 6377 9333 6411 9367
rect 8033 9333 8067 9367
rect 8217 9333 8251 9367
rect 8953 9333 8987 9367
rect 10149 9333 10183 9367
rect 10425 9333 10459 9367
rect 3065 9129 3099 9163
rect 7849 9129 7883 9163
rect 9229 9129 9263 9163
rect 10057 9129 10091 9163
rect 9781 8993 9815 9027
rect 4169 8925 4203 8959
rect 4445 8925 4479 8959
rect 6009 8925 6043 8959
rect 7757 8925 7791 8959
rect 8033 8925 8067 8959
rect 8217 8925 8251 8959
rect 9597 8925 9631 8959
rect 2697 8857 2731 8891
rect 2881 8857 2915 8891
rect 4261 8857 4295 8891
rect 6254 8857 6288 8891
rect 9413 8857 9447 8891
rect 10241 8857 10275 8891
rect 4629 8789 4663 8823
rect 7389 8789 7423 8823
rect 7573 8789 7607 8823
rect 8401 8789 8435 8823
rect 9505 8789 9539 8823
rect 9873 8789 9907 8823
rect 10041 8789 10075 8823
rect 2789 8585 2823 8619
rect 4829 8585 4863 8619
rect 8401 8585 8435 8619
rect 10031 8585 10065 8619
rect 4629 8517 4663 8551
rect 10241 8517 10275 8551
rect 1409 8449 1443 8483
rect 1676 8449 1710 8483
rect 5733 8449 5767 8483
rect 9525 8449 9559 8483
rect 9781 8381 9815 8415
rect 9873 8313 9907 8347
rect 4813 8245 4847 8279
rect 4997 8245 5031 8279
rect 5549 8245 5583 8279
rect 10057 8245 10091 8279
rect 5549 8041 5583 8075
rect 3893 7973 3927 8007
rect 5017 7837 5051 7871
rect 5273 7837 5307 7871
rect 5917 7837 5951 7871
rect 9137 7815 9171 7849
rect 9413 7837 9447 7871
rect 10241 7837 10275 7871
rect 5549 7769 5583 7803
rect 9597 7769 9631 7803
rect 5365 7701 5399 7735
rect 9229 7701 9263 7735
rect 10425 7701 10459 7735
rect 2697 7497 2731 7531
rect 6561 7497 6595 7531
rect 9781 7497 9815 7531
rect 4988 7429 5022 7463
rect 9965 7429 9999 7463
rect 1501 7361 1535 7395
rect 3821 7361 3855 7395
rect 4629 7361 4663 7395
rect 6377 7361 6411 7395
rect 7941 7361 7975 7395
rect 4077 7293 4111 7327
rect 4721 7293 4755 7327
rect 6101 7225 6135 7259
rect 10333 7225 10367 7259
rect 1593 7157 1627 7191
rect 4537 7157 4571 7191
rect 9229 7157 9263 7191
rect 9965 7157 9999 7191
rect 3433 6953 3467 6987
rect 3801 6953 3835 6987
rect 6929 6953 6963 6987
rect 2329 6817 2363 6851
rect 1777 6749 1811 6783
rect 1961 6749 1995 6783
rect 2053 6749 2087 6783
rect 2145 6749 2179 6783
rect 2605 6749 2639 6783
rect 2881 6749 2915 6783
rect 5181 6749 5215 6783
rect 8401 6749 8435 6783
rect 9505 6749 9539 6783
rect 9689 6749 9723 6783
rect 10241 6749 10275 6783
rect 3249 6681 3283 6715
rect 4936 6681 4970 6715
rect 5641 6681 5675 6715
rect 1593 6613 1627 6647
rect 2329 6613 2363 6647
rect 2421 6613 2455 6647
rect 2789 6613 2823 6647
rect 3449 6613 3483 6647
rect 3617 6613 3651 6647
rect 8217 6613 8251 6647
rect 9597 6613 9631 6647
rect 10425 6613 10459 6647
rect 1685 6409 1719 6443
rect 1961 6409 1995 6443
rect 6469 6409 6503 6443
rect 8493 6409 8527 6443
rect 8861 6409 8895 6443
rect 8953 6409 8987 6443
rect 10057 6409 10091 6443
rect 2697 6341 2731 6375
rect 2913 6341 2947 6375
rect 5733 6341 5767 6375
rect 6009 6341 6043 6375
rect 6193 6341 6227 6375
rect 7380 6341 7414 6375
rect 8585 6341 8619 6375
rect 9381 6341 9415 6375
rect 9597 6341 9631 6375
rect 9689 6341 9723 6375
rect 9873 6341 9907 6375
rect 1501 6273 1535 6307
rect 1777 6273 1811 6307
rect 1961 6273 1995 6307
rect 3157 6273 3191 6307
rect 3341 6273 3375 6307
rect 3433 6273 3467 6307
rect 3525 6273 3559 6307
rect 3709 6273 3743 6307
rect 5917 6273 5951 6307
rect 6653 6273 6687 6307
rect 8769 6273 8803 6307
rect 3985 6205 4019 6239
rect 6837 6205 6871 6239
rect 7113 6205 7147 6239
rect 5917 6137 5951 6171
rect 2881 6069 2915 6103
rect 3065 6069 3099 6103
rect 3893 6069 3927 6103
rect 9137 6069 9171 6103
rect 9229 6069 9263 6103
rect 9413 6069 9447 6103
rect 1501 5865 1535 5899
rect 4721 5865 4755 5899
rect 6101 5865 6135 5899
rect 7389 5865 7423 5899
rect 6285 5797 6319 5831
rect 9413 5797 9447 5831
rect 9505 5797 9539 5831
rect 2881 5729 2915 5763
rect 2625 5661 2659 5695
rect 4905 5661 4939 5695
rect 5089 5661 5123 5695
rect 5273 5661 5307 5695
rect 5365 5661 5399 5695
rect 5457 5661 5491 5695
rect 6377 5661 6411 5695
rect 6653 5661 6687 5695
rect 6929 5661 6963 5695
rect 7113 5661 7147 5695
rect 8769 5661 8803 5695
rect 9137 5661 9171 5695
rect 9689 5661 9723 5695
rect 10241 5661 10275 5695
rect 5917 5593 5951 5627
rect 6837 5593 6871 5627
rect 8502 5593 8536 5627
rect 9413 5593 9447 5627
rect 5733 5525 5767 5559
rect 6117 5525 6151 5559
rect 6469 5525 6503 5559
rect 6929 5525 6963 5559
rect 9229 5525 9263 5559
rect 10425 5525 10459 5559
rect 1961 5321 1995 5355
rect 5549 5321 5583 5355
rect 5733 5321 5767 5355
rect 5901 5321 5935 5355
rect 10123 5321 10157 5355
rect 1777 5253 1811 5287
rect 2881 5253 2915 5287
rect 6101 5253 6135 5287
rect 10333 5253 10367 5287
rect 1409 5185 1443 5219
rect 2697 5185 2731 5219
rect 4914 5185 4948 5219
rect 5457 5185 5491 5219
rect 5641 5185 5675 5219
rect 7674 5185 7708 5219
rect 8217 5185 8251 5219
rect 9422 5185 9456 5219
rect 9689 5185 9723 5219
rect 3065 5117 3099 5151
rect 5181 5117 5215 5151
rect 7941 5117 7975 5151
rect 8033 5049 8067 5083
rect 1777 4981 1811 5015
rect 3801 4981 3835 5015
rect 5917 4981 5951 5015
rect 6561 4981 6595 5015
rect 8309 4981 8343 5015
rect 9965 4981 9999 5015
rect 10149 4981 10183 5015
rect 2881 4777 2915 4811
rect 3065 4777 3099 4811
rect 4353 4777 4387 4811
rect 5089 4777 5123 4811
rect 5273 4777 5307 4811
rect 6285 4777 6319 4811
rect 8033 4777 8067 4811
rect 3525 4641 3559 4675
rect 2605 4573 2639 4607
rect 3341 4573 3375 4607
rect 4261 4573 4295 4607
rect 4445 4573 4479 4607
rect 6101 4573 6135 4607
rect 6377 4573 6411 4607
rect 6653 4573 6687 4607
rect 10241 4573 10275 4607
rect 4905 4505 4939 4539
rect 5105 4505 5139 4539
rect 6898 4505 6932 4539
rect 3157 4437 3191 4471
rect 6561 4437 6595 4471
rect 10425 4437 10459 4471
rect 2230 4233 2264 4267
rect 2789 4233 2823 4267
rect 1593 4165 1627 4199
rect 2421 4165 2455 4199
rect 2605 4165 2639 4199
rect 6837 4165 6871 4199
rect 7037 4165 7071 4199
rect 7633 4165 7667 4199
rect 7849 4165 7883 4199
rect 1777 4097 1811 4131
rect 2053 4097 2087 4131
rect 2145 4097 2179 4131
rect 2329 4097 2363 4131
rect 2697 4097 2731 4131
rect 4997 4097 5031 4131
rect 4813 4029 4847 4063
rect 5089 4029 5123 4063
rect 5181 4029 5215 4063
rect 5273 4029 5307 4063
rect 1961 3961 1995 3995
rect 7205 3961 7239 3995
rect 2973 3893 3007 3927
rect 7021 3893 7055 3927
rect 7481 3893 7515 3927
rect 7665 3893 7699 3927
rect 4813 3689 4847 3723
rect 7021 3689 7055 3723
rect 9873 3689 9907 3723
rect 7205 3621 7239 3655
rect 7389 3621 7423 3655
rect 9321 3621 9355 3655
rect 2053 3553 2087 3587
rect 5641 3553 5675 3587
rect 7665 3553 7699 3587
rect 2145 3485 2179 3519
rect 2973 3485 3007 3519
rect 4721 3485 4755 3519
rect 4997 3485 5031 3519
rect 5181 3485 5215 3519
rect 5549 3485 5583 3519
rect 5897 3485 5931 3519
rect 9045 3485 9079 3519
rect 9505 3485 9539 3519
rect 10241 3485 10275 3519
rect 9321 3417 9355 3451
rect 9689 3417 9723 3451
rect 3157 3349 3191 3383
rect 9137 3349 9171 3383
rect 10425 3349 10459 3383
rect 2789 3145 2823 3179
rect 4261 3145 4295 3179
rect 5733 3145 5767 3179
rect 6561 3145 6595 3179
rect 8401 3145 8435 3179
rect 9413 3145 9447 3179
rect 4620 3077 4654 3111
rect 1409 3009 1443 3043
rect 1676 3009 1710 3043
rect 3065 3009 3099 3043
rect 3249 3009 3283 3043
rect 3893 3009 3927 3043
rect 4077 3009 4111 3043
rect 6377 3009 6411 3043
rect 7021 3009 7055 3043
rect 7277 3009 7311 3043
rect 9413 3009 9447 3043
rect 9781 3009 9815 3043
rect 10057 3009 10091 3043
rect 10149 3009 10183 3043
rect 10333 3009 10367 3043
rect 4353 2941 4387 2975
rect 2881 2805 2915 2839
rect 2421 2601 2455 2635
rect 5365 2601 5399 2635
rect 2513 2533 2547 2567
rect 4997 2533 5031 2567
rect 6101 2533 6135 2567
rect 2145 2465 2179 2499
rect 2237 2465 2271 2499
rect 1961 2397 1995 2431
rect 2053 2397 2087 2431
rect 2513 2397 2547 2431
rect 2697 2397 2731 2431
rect 5917 2397 5951 2431
rect 6101 2397 6135 2431
rect 9965 2397 9999 2431
rect 10241 2397 10275 2431
rect 5365 2329 5399 2363
rect 5549 2261 5583 2295
rect 10149 2261 10183 2295
rect 10425 2261 10459 2295
<< metal1 >>
rect 1670 11568 1676 11620
rect 1728 11608 1734 11620
rect 8570 11608 8576 11620
rect 1728 11580 8576 11608
rect 1728 11568 1734 11580
rect 8570 11568 8576 11580
rect 8628 11568 8634 11620
rect 2590 11500 2596 11552
rect 2648 11540 2654 11552
rect 4522 11540 4528 11552
rect 2648 11512 4528 11540
rect 2648 11500 2654 11512
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 1104 11450 10764 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 6950 11450
rect 7002 11398 7014 11450
rect 7066 11398 7078 11450
rect 7130 11398 7142 11450
rect 7194 11398 7206 11450
rect 7258 11398 10764 11450
rect 1104 11376 10764 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 1670 11336 1676 11348
rect 1627 11308 1676 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 3476 11308 4077 11336
rect 3476 11296 3482 11308
rect 4065 11305 4077 11308
rect 4111 11305 4123 11339
rect 4065 11299 4123 11305
rect 4172 11308 4476 11336
rect 1762 11228 1768 11280
rect 1820 11268 1826 11280
rect 3050 11268 3056 11280
rect 1820 11240 3056 11268
rect 1820 11228 1826 11240
rect 1578 11160 1584 11212
rect 1636 11200 1642 11212
rect 2409 11203 2467 11209
rect 2409 11200 2421 11203
rect 1636 11172 2421 11200
rect 1636 11160 1642 11172
rect 2409 11169 2421 11172
rect 2455 11169 2467 11203
rect 2409 11163 2467 11169
rect 2590 11160 2596 11212
rect 2648 11160 2654 11212
rect 2700 11209 2728 11240
rect 3050 11228 3056 11240
rect 3108 11228 3114 11280
rect 3142 11228 3148 11280
rect 3200 11268 3206 11280
rect 3329 11271 3387 11277
rect 3329 11268 3341 11271
rect 3200 11240 3341 11268
rect 3200 11228 3206 11240
rect 3329 11237 3341 11240
rect 3375 11237 3387 11271
rect 3329 11231 3387 11237
rect 3694 11228 3700 11280
rect 3752 11268 3758 11280
rect 4172 11268 4200 11308
rect 3752 11240 4200 11268
rect 3752 11228 3758 11240
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11169 2743 11203
rect 2685 11163 2743 11169
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 4154 11200 4160 11212
rect 2823 11172 4160 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 1486 11092 1492 11144
rect 1544 11092 1550 11144
rect 1854 11092 1860 11144
rect 1912 11132 1918 11144
rect 2608 11132 2636 11160
rect 1912 11104 2636 11132
rect 1912 11092 1918 11104
rect 2498 11024 2504 11076
rect 2556 11064 2562 11076
rect 2792 11064 2820 11163
rect 4154 11160 4160 11172
rect 4212 11160 4218 11212
rect 4448 11200 4476 11308
rect 8478 11296 8484 11348
rect 8536 11296 8542 11348
rect 9674 11336 9680 11348
rect 8588 11308 9680 11336
rect 5261 11271 5319 11277
rect 5261 11237 5273 11271
rect 5307 11268 5319 11271
rect 5626 11268 5632 11280
rect 5307 11240 5632 11268
rect 5307 11237 5319 11240
rect 5261 11231 5319 11237
rect 5626 11228 5632 11240
rect 5684 11228 5690 11280
rect 8386 11268 8392 11280
rect 5736 11240 8392 11268
rect 5736 11200 5764 11240
rect 8386 11228 8392 11240
rect 8444 11228 8450 11280
rect 8588 11200 8616 11308
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 8754 11228 8760 11280
rect 8812 11228 8818 11280
rect 4448 11172 5764 11200
rect 8312 11172 8616 11200
rect 4448 11141 4476 11172
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11132 2927 11135
rect 4341 11135 4399 11141
rect 2915 11104 3832 11132
rect 2915 11101 2927 11104
rect 2869 11095 2927 11101
rect 3804 11076 3832 11104
rect 4341 11101 4353 11135
rect 4387 11101 4399 11135
rect 4341 11095 4399 11101
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 2556 11036 2820 11064
rect 2556 11024 2562 11036
rect 3050 11024 3056 11076
rect 3108 11064 3114 11076
rect 3694 11064 3700 11076
rect 3108 11036 3700 11064
rect 3108 11024 3114 11036
rect 3694 11024 3700 11036
rect 3752 11024 3758 11076
rect 3786 11024 3792 11076
rect 3844 11064 3850 11076
rect 4356 11064 4384 11095
rect 5718 11092 5724 11144
rect 5776 11092 5782 11144
rect 5810 11092 5816 11144
rect 5868 11092 5874 11144
rect 8312 11141 8340 11172
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 8573 11135 8631 11141
rect 8573 11132 8585 11135
rect 8536 11104 8585 11132
rect 8536 11092 8542 11104
rect 8573 11101 8585 11104
rect 8619 11101 8631 11135
rect 8573 11095 8631 11101
rect 8941 11135 8999 11141
rect 8941 11101 8953 11135
rect 8987 11132 8999 11135
rect 8987 11104 9444 11132
rect 8987 11101 8999 11104
rect 8941 11095 8999 11101
rect 9416 11076 9444 11104
rect 3844 11036 4384 11064
rect 3844 11024 3850 11036
rect 4614 11024 4620 11076
rect 4672 11024 4678 11076
rect 5534 11024 5540 11076
rect 5592 11024 5598 11076
rect 7466 11024 7472 11076
rect 7524 11064 7530 11076
rect 9186 11067 9244 11073
rect 9186 11064 9198 11067
rect 7524 11036 9198 11064
rect 7524 11024 7530 11036
rect 9186 11033 9198 11036
rect 9232 11033 9244 11067
rect 9186 11027 9244 11033
rect 9398 11024 9404 11076
rect 9456 11024 9462 11076
rect 3510 10956 3516 11008
rect 3568 10956 3574 11008
rect 4249 10999 4307 11005
rect 4249 10965 4261 10999
rect 4295 10996 4307 10999
rect 4522 10996 4528 11008
rect 4295 10968 4528 10996
rect 4295 10965 4307 10968
rect 4249 10959 4307 10965
rect 4522 10956 4528 10968
rect 4580 10996 4586 11008
rect 5718 10996 5724 11008
rect 4580 10968 5724 10996
rect 4580 10956 4586 10968
rect 5718 10956 5724 10968
rect 5776 10956 5782 11008
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 10042 10996 10048 11008
rect 7248 10968 10048 10996
rect 7248 10956 7254 10968
rect 10042 10956 10048 10968
rect 10100 10996 10106 11008
rect 10321 10999 10379 11005
rect 10321 10996 10333 10999
rect 10100 10968 10333 10996
rect 10100 10956 10106 10968
rect 10321 10965 10333 10968
rect 10367 10965 10379 10999
rect 10321 10959 10379 10965
rect 1104 10906 10764 10928
rect 1104 10854 2610 10906
rect 2662 10854 2674 10906
rect 2726 10854 2738 10906
rect 2790 10854 2802 10906
rect 2854 10854 2866 10906
rect 2918 10854 7610 10906
rect 7662 10854 7674 10906
rect 7726 10854 7738 10906
rect 7790 10854 7802 10906
rect 7854 10854 7866 10906
rect 7918 10854 10764 10906
rect 1104 10832 10764 10854
rect 1762 10752 1768 10804
rect 1820 10752 1826 10804
rect 1854 10752 1860 10804
rect 1912 10752 1918 10804
rect 3142 10792 3148 10804
rect 2700 10764 3148 10792
rect 1780 10724 1808 10752
rect 2700 10733 2728 10764
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 7190 10792 7196 10804
rect 4120 10764 7196 10792
rect 4120 10752 4126 10764
rect 7190 10752 7196 10764
rect 7248 10752 7254 10804
rect 7377 10795 7435 10801
rect 7377 10761 7389 10795
rect 7423 10792 7435 10795
rect 7926 10792 7932 10804
rect 7423 10764 7932 10792
rect 7423 10761 7435 10764
rect 7377 10755 7435 10761
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 8021 10795 8079 10801
rect 8021 10761 8033 10795
rect 8067 10761 8079 10795
rect 8021 10755 8079 10761
rect 8481 10795 8539 10801
rect 8481 10761 8493 10795
rect 8527 10792 8539 10795
rect 9582 10792 9588 10804
rect 8527 10764 9588 10792
rect 8527 10761 8539 10764
rect 8481 10755 8539 10761
rect 2469 10727 2527 10733
rect 2469 10724 2481 10727
rect 1780 10696 2481 10724
rect 2469 10693 2481 10696
rect 2515 10693 2527 10727
rect 2469 10687 2527 10693
rect 2685 10727 2743 10733
rect 2685 10693 2697 10727
rect 2731 10693 2743 10727
rect 2685 10687 2743 10693
rect 2884 10696 3280 10724
rect 1486 10616 1492 10668
rect 1544 10656 1550 10668
rect 1670 10656 1676 10668
rect 1544 10628 1676 10656
rect 1544 10616 1550 10628
rect 1670 10616 1676 10628
rect 1728 10616 1734 10668
rect 2884 10665 2912 10696
rect 3252 10668 3280 10696
rect 4154 10684 4160 10736
rect 4212 10724 4218 10736
rect 4614 10724 4620 10736
rect 4212 10696 4620 10724
rect 4212 10684 4218 10696
rect 4614 10684 4620 10696
rect 4672 10724 4678 10736
rect 5626 10724 5632 10736
rect 4672 10696 5632 10724
rect 4672 10684 4678 10696
rect 5626 10684 5632 10696
rect 5684 10724 5690 10736
rect 8036 10724 8064 10755
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 9278 10727 9336 10733
rect 9278 10724 9290 10727
rect 5684 10696 7972 10724
rect 8036 10696 9290 10724
rect 5684 10684 5690 10696
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 2869 10659 2927 10665
rect 1811 10628 2820 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 1974 10591 2032 10597
rect 1974 10557 1986 10591
rect 2020 10588 2032 10591
rect 2498 10588 2504 10600
rect 2020 10560 2504 10588
rect 2020 10557 2032 10560
rect 1974 10551 2032 10557
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 2792 10588 2820 10628
rect 2869 10625 2881 10659
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 3050 10616 3056 10668
rect 3108 10616 3114 10668
rect 3234 10616 3240 10668
rect 3292 10616 3298 10668
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 5810 10656 5816 10668
rect 3936 10628 5816 10656
rect 3936 10616 3942 10628
rect 5810 10616 5816 10628
rect 5868 10616 5874 10668
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 7650 10656 7656 10668
rect 7515 10628 7656 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 7834 10616 7840 10668
rect 7892 10616 7898 10668
rect 7944 10656 7972 10696
rect 9278 10693 9290 10696
rect 9324 10693 9336 10727
rect 9278 10687 9336 10693
rect 9398 10684 9404 10736
rect 9456 10684 9462 10736
rect 7944 10628 8156 10656
rect 3786 10588 3792 10600
rect 2792 10560 3792 10588
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 7101 10591 7159 10597
rect 7101 10557 7113 10591
rect 7147 10557 7159 10591
rect 7101 10551 7159 10557
rect 7561 10591 7619 10597
rect 7561 10557 7573 10591
rect 7607 10588 7619 10591
rect 8018 10588 8024 10600
rect 7607 10560 8024 10588
rect 7607 10557 7619 10560
rect 7561 10551 7619 10557
rect 5994 10520 6000 10532
rect 2746 10492 6000 10520
rect 1854 10412 1860 10464
rect 1912 10452 1918 10464
rect 2133 10455 2191 10461
rect 2133 10452 2145 10455
rect 1912 10424 2145 10452
rect 1912 10412 1918 10424
rect 2133 10421 2145 10424
rect 2179 10421 2191 10455
rect 2133 10415 2191 10421
rect 2314 10412 2320 10464
rect 2372 10412 2378 10464
rect 2501 10455 2559 10461
rect 2501 10421 2513 10455
rect 2547 10452 2559 10455
rect 2746 10452 2774 10492
rect 5994 10480 6000 10492
rect 6052 10480 6058 10532
rect 6362 10480 6368 10532
rect 6420 10520 6426 10532
rect 7116 10520 7144 10551
rect 8018 10548 8024 10560
rect 8076 10548 8082 10600
rect 8128 10588 8156 10628
rect 8294 10616 8300 10668
rect 8352 10616 8358 10668
rect 8386 10616 8392 10668
rect 8444 10656 8450 10668
rect 8573 10659 8631 10665
rect 8573 10656 8585 10659
rect 8444 10628 8585 10656
rect 8444 10616 8450 10628
rect 8573 10625 8585 10628
rect 8619 10656 8631 10659
rect 8662 10656 8668 10668
rect 8619 10628 8668 10656
rect 8619 10625 8631 10628
rect 8573 10619 8631 10625
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 8757 10659 8815 10665
rect 8757 10625 8769 10659
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 9033 10659 9091 10665
rect 9033 10625 9045 10659
rect 9079 10656 9091 10659
rect 9416 10656 9444 10684
rect 9079 10628 9444 10656
rect 9079 10625 9091 10628
rect 9033 10619 9091 10625
rect 8772 10588 8800 10619
rect 8128 10560 8800 10588
rect 8202 10520 8208 10532
rect 6420 10492 8208 10520
rect 6420 10480 6426 10492
rect 8202 10480 8208 10492
rect 8260 10480 8266 10532
rect 8478 10480 8484 10532
rect 8536 10520 8542 10532
rect 8536 10492 9076 10520
rect 8536 10480 8542 10492
rect 2547 10424 2774 10452
rect 2961 10455 3019 10461
rect 2547 10421 2559 10424
rect 2501 10415 2559 10421
rect 2961 10421 2973 10455
rect 3007 10452 3019 10455
rect 3510 10452 3516 10464
rect 3007 10424 3516 10452
rect 3007 10421 3019 10424
rect 2961 10415 3019 10421
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 3694 10412 3700 10464
rect 3752 10452 3758 10464
rect 6454 10452 6460 10464
rect 3752 10424 6460 10452
rect 3752 10412 3758 10424
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 7745 10455 7803 10461
rect 7745 10421 7757 10455
rect 7791 10452 7803 10455
rect 8846 10452 8852 10464
rect 7791 10424 8852 10452
rect 7791 10421 7803 10424
rect 7745 10415 7803 10421
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 8938 10412 8944 10464
rect 8996 10412 9002 10464
rect 9048 10452 9076 10492
rect 10413 10455 10471 10461
rect 10413 10452 10425 10455
rect 9048 10424 10425 10452
rect 10413 10421 10425 10424
rect 10459 10421 10471 10455
rect 10413 10415 10471 10421
rect 1104 10362 10764 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 6950 10362
rect 7002 10310 7014 10362
rect 7066 10310 7078 10362
rect 7130 10310 7142 10362
rect 7194 10310 7206 10362
rect 7258 10310 10764 10362
rect 1104 10288 10764 10310
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 3970 10248 3976 10260
rect 2924 10220 3976 10248
rect 2924 10208 2930 10220
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 4522 10208 4528 10260
rect 4580 10208 4586 10260
rect 4709 10251 4767 10257
rect 4709 10217 4721 10251
rect 4755 10248 4767 10251
rect 7834 10248 7840 10260
rect 4755 10220 7840 10248
rect 4755 10217 4767 10220
rect 4709 10211 4767 10217
rect 7834 10208 7840 10220
rect 7892 10208 7898 10260
rect 7926 10208 7932 10260
rect 7984 10248 7990 10260
rect 8478 10248 8484 10260
rect 7984 10220 8484 10248
rect 7984 10208 7990 10220
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 9217 10251 9275 10257
rect 9217 10248 9229 10251
rect 8628 10220 9229 10248
rect 8628 10208 8634 10220
rect 9217 10217 9229 10220
rect 9263 10248 9275 10251
rect 9858 10248 9864 10260
rect 9263 10220 9864 10248
rect 9263 10217 9275 10220
rect 9217 10211 9275 10217
rect 9858 10208 9864 10220
rect 9916 10248 9922 10260
rect 10870 10248 10876 10260
rect 9916 10220 10876 10248
rect 9916 10208 9922 10220
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 3145 10183 3203 10189
rect 3145 10149 3157 10183
rect 3191 10180 3203 10183
rect 6270 10180 6276 10192
rect 3191 10152 6276 10180
rect 3191 10149 3203 10152
rect 3145 10143 3203 10149
rect 6270 10140 6276 10152
rect 6328 10140 6334 10192
rect 9140 10152 9674 10180
rect 2593 10115 2651 10121
rect 2593 10081 2605 10115
rect 2639 10112 2651 10115
rect 2639 10084 3188 10112
rect 2639 10081 2651 10084
rect 2593 10075 2651 10081
rect 3160 10056 3188 10084
rect 3602 10072 3608 10124
rect 3660 10072 3666 10124
rect 3896 10084 5028 10112
rect 1670 10004 1676 10056
rect 1728 10004 1734 10056
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10044 2927 10047
rect 2958 10044 2964 10056
rect 2915 10016 2964 10044
rect 2915 10013 2927 10016
rect 2869 10007 2927 10013
rect 2958 10004 2964 10016
rect 3016 10004 3022 10056
rect 3142 10004 3148 10056
rect 3200 10004 3206 10056
rect 3418 10004 3424 10056
rect 3476 10004 3482 10056
rect 3694 10004 3700 10056
rect 3752 10044 3758 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3752 10016 3801 10044
rect 3752 10004 3758 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 934 9936 940 9988
rect 992 9976 998 9988
rect 3896 9976 3924 10084
rect 4062 10004 4068 10056
rect 4120 10004 4126 10056
rect 4614 10004 4620 10056
rect 4672 10004 4678 10056
rect 4798 10004 4804 10056
rect 4856 10004 4862 10056
rect 5000 10053 5028 10084
rect 6086 10072 6092 10124
rect 6144 10112 6150 10124
rect 6144 10084 6316 10112
rect 6144 10072 6150 10084
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10044 6055 10047
rect 6178 10044 6184 10056
rect 6043 10016 6184 10044
rect 6043 10013 6055 10016
rect 5997 10007 6055 10013
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6288 10053 6316 10084
rect 7650 10072 7656 10124
rect 7708 10112 7714 10124
rect 8294 10112 8300 10124
rect 7708 10084 8300 10112
rect 7708 10072 7714 10084
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 8573 10115 8631 10121
rect 8573 10081 8585 10115
rect 8619 10112 8631 10115
rect 9140 10112 9168 10152
rect 8619 10084 9168 10112
rect 9646 10112 9674 10152
rect 9646 10084 10272 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 6638 10044 6644 10056
rect 6595 10016 6644 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 6638 10004 6644 10016
rect 6696 10004 6702 10056
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 9030 10044 9036 10056
rect 8076 10016 9036 10044
rect 8076 10004 8082 10016
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 9122 10004 9128 10056
rect 9180 10044 9186 10056
rect 9180 10016 9996 10044
rect 9180 10004 9186 10016
rect 992 9948 3924 9976
rect 4341 9979 4399 9985
rect 992 9936 998 9948
rect 4341 9945 4353 9979
rect 4387 9976 4399 9979
rect 4632 9976 4660 10004
rect 4387 9948 4660 9976
rect 4387 9945 4399 9948
rect 4341 9939 4399 9945
rect 4706 9936 4712 9988
rect 4764 9976 4770 9988
rect 6794 9979 6852 9985
rect 6794 9976 6806 9979
rect 4764 9948 6806 9976
rect 4764 9936 4770 9948
rect 6794 9945 6806 9948
rect 6840 9945 6852 9979
rect 6794 9939 6852 9945
rect 6914 9936 6920 9988
rect 6972 9976 6978 9988
rect 9766 9976 9772 9988
rect 6972 9948 9772 9976
rect 6972 9936 6978 9948
rect 1489 9911 1547 9917
rect 1489 9877 1501 9911
rect 1535 9908 1547 9911
rect 1670 9908 1676 9920
rect 1535 9880 1676 9908
rect 1535 9877 1547 9880
rect 1489 9871 1547 9877
rect 1670 9868 1676 9880
rect 1728 9868 1734 9920
rect 2498 9868 2504 9920
rect 2556 9908 2562 9920
rect 2777 9911 2835 9917
rect 2777 9908 2789 9911
rect 2556 9880 2789 9908
rect 2556 9868 2562 9880
rect 2777 9877 2789 9880
rect 2823 9877 2835 9911
rect 2777 9871 2835 9877
rect 2866 9868 2872 9920
rect 2924 9908 2930 9920
rect 2961 9911 3019 9917
rect 2961 9908 2973 9911
rect 2924 9880 2973 9908
rect 2924 9868 2930 9880
rect 2961 9877 2973 9880
rect 3007 9877 3019 9911
rect 2961 9871 3019 9877
rect 3234 9868 3240 9920
rect 3292 9868 3298 9920
rect 3326 9868 3332 9920
rect 3384 9908 3390 9920
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 3384 9880 3893 9908
rect 3384 9868 3390 9880
rect 3881 9877 3893 9880
rect 3927 9877 3939 9911
rect 3881 9871 3939 9877
rect 4246 9868 4252 9920
rect 4304 9868 4310 9920
rect 4430 9868 4436 9920
rect 4488 9908 4494 9920
rect 4541 9911 4599 9917
rect 4541 9908 4553 9911
rect 4488 9880 4553 9908
rect 4488 9868 4494 9880
rect 4541 9877 4553 9880
rect 4587 9877 4599 9911
rect 4541 9871 4599 9877
rect 4890 9868 4896 9920
rect 4948 9868 4954 9920
rect 6086 9868 6092 9920
rect 6144 9868 6150 9920
rect 6457 9911 6515 9917
rect 6457 9877 6469 9911
rect 6503 9908 6515 9911
rect 7374 9908 7380 9920
rect 6503 9880 7380 9908
rect 6503 9877 6515 9880
rect 6457 9871 6515 9877
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 7944 9917 7972 9948
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 9858 9936 9864 9988
rect 9916 9936 9922 9988
rect 9968 9985 9996 10016
rect 10244 9985 10272 10084
rect 9953 9979 10011 9985
rect 9953 9945 9965 9979
rect 9999 9945 10011 9979
rect 9953 9939 10011 9945
rect 10229 9979 10287 9985
rect 10229 9945 10241 9979
rect 10275 9976 10287 9979
rect 10275 9948 10824 9976
rect 10275 9945 10287 9948
rect 10229 9939 10287 9945
rect 10796 9920 10824 9948
rect 7929 9911 7987 9917
rect 7929 9877 7941 9911
rect 7975 9877 7987 9911
rect 7929 9871 7987 9877
rect 8294 9868 8300 9920
rect 8352 9908 8358 9920
rect 9214 9908 9220 9920
rect 8352 9880 9220 9908
rect 8352 9868 8358 9880
rect 9214 9868 9220 9880
rect 9272 9868 9278 9920
rect 9582 9868 9588 9920
rect 9640 9908 9646 9920
rect 9677 9911 9735 9917
rect 9677 9908 9689 9911
rect 9640 9880 9689 9908
rect 9640 9868 9646 9880
rect 9677 9877 9689 9880
rect 9723 9877 9735 9911
rect 9677 9871 9735 9877
rect 10045 9911 10103 9917
rect 10045 9877 10057 9911
rect 10091 9908 10103 9911
rect 10686 9908 10692 9920
rect 10091 9880 10692 9908
rect 10091 9877 10103 9880
rect 10045 9871 10103 9877
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 10778 9868 10784 9920
rect 10836 9868 10842 9920
rect 1104 9818 10764 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 7610 9818
rect 7662 9766 7674 9818
rect 7726 9766 7738 9818
rect 7790 9766 7802 9818
rect 7854 9766 7866 9818
rect 7918 9766 10764 9818
rect 1104 9744 10764 9766
rect 2501 9707 2559 9713
rect 2501 9673 2513 9707
rect 2547 9704 2559 9707
rect 4706 9704 4712 9716
rect 2547 9676 4712 9704
rect 2547 9673 2559 9676
rect 2501 9667 2559 9673
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 5994 9664 6000 9716
rect 6052 9664 6058 9716
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 8018 9704 8024 9716
rect 7616 9676 8024 9704
rect 7616 9664 7622 9676
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 8220 9676 9076 9704
rect 3237 9639 3295 9645
rect 3237 9605 3249 9639
rect 3283 9636 3295 9639
rect 4614 9636 4620 9648
rect 3283 9608 4620 9636
rect 3283 9605 3295 9608
rect 3237 9599 3295 9605
rect 4614 9596 4620 9608
rect 4672 9596 4678 9648
rect 4890 9596 4896 9648
rect 4948 9645 4954 9648
rect 4948 9636 4960 9645
rect 4948 9608 4993 9636
rect 4948 9599 4960 9608
rect 4948 9596 4954 9599
rect 6638 9596 6644 9648
rect 6696 9636 6702 9648
rect 8220 9645 8248 9676
rect 8205 9639 8263 9645
rect 6696 9608 7788 9636
rect 6696 9596 6702 9608
rect 658 9528 664 9580
rect 716 9568 722 9580
rect 1857 9571 1915 9577
rect 1857 9568 1869 9571
rect 716 9540 1869 9568
rect 716 9528 722 9540
rect 1857 9537 1869 9540
rect 1903 9537 1915 9571
rect 1857 9531 1915 9537
rect 2314 9528 2320 9580
rect 2372 9528 2378 9580
rect 4430 9568 4436 9580
rect 3436 9540 4436 9568
rect 3436 9441 3464 9540
rect 4430 9528 4436 9540
rect 4488 9528 4494 9580
rect 5074 9528 5080 9580
rect 5132 9568 5138 9580
rect 5997 9571 6055 9577
rect 5997 9568 6009 9571
rect 5132 9540 6009 9568
rect 5132 9528 5138 9540
rect 5997 9537 6009 9540
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9537 6239 9571
rect 6914 9568 6920 9580
rect 6181 9531 6239 9537
rect 6380 9540 6920 9568
rect 3694 9460 3700 9512
rect 3752 9500 3758 9512
rect 4062 9500 4068 9512
rect 3752 9472 4068 9500
rect 3752 9460 3758 9472
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 5169 9503 5227 9509
rect 5169 9469 5181 9503
rect 5215 9469 5227 9503
rect 6196 9500 6224 9531
rect 5169 9463 5227 9469
rect 5828 9472 6224 9500
rect 2869 9435 2927 9441
rect 2869 9401 2881 9435
rect 2915 9432 2927 9435
rect 3421 9435 3479 9441
rect 2915 9404 3004 9432
rect 2915 9401 2927 9404
rect 2869 9395 2927 9401
rect 2976 9376 3004 9404
rect 3421 9401 3433 9435
rect 3467 9401 3479 9435
rect 4154 9432 4160 9444
rect 3421 9395 3479 9401
rect 3712 9404 4160 9432
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 2774 9364 2780 9376
rect 2087 9336 2780 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 2774 9324 2780 9336
rect 2832 9324 2838 9376
rect 2958 9324 2964 9376
rect 3016 9324 3022 9376
rect 3237 9367 3295 9373
rect 3237 9333 3249 9367
rect 3283 9364 3295 9367
rect 3712 9364 3740 9404
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 3283 9336 3740 9364
rect 3789 9367 3847 9373
rect 3283 9333 3295 9336
rect 3237 9327 3295 9333
rect 3789 9333 3801 9367
rect 3835 9364 3847 9367
rect 3970 9364 3976 9376
rect 3835 9336 3976 9364
rect 3835 9333 3847 9336
rect 3789 9327 3847 9333
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 5184 9364 5212 9463
rect 5828 9376 5856 9472
rect 5994 9392 6000 9444
rect 6052 9432 6058 9444
rect 6380 9432 6408 9540
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7489 9571 7547 9577
rect 7489 9537 7501 9571
rect 7535 9568 7547 9571
rect 7650 9568 7656 9580
rect 7535 9540 7656 9568
rect 7535 9537 7547 9540
rect 7489 9531 7547 9537
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7760 9509 7788 9608
rect 8205 9605 8217 9639
rect 8251 9605 8263 9639
rect 8205 9599 8263 9605
rect 8294 9596 8300 9648
rect 8352 9636 8358 9648
rect 8941 9639 8999 9645
rect 8941 9636 8953 9639
rect 8352 9608 8953 9636
rect 8352 9596 8358 9608
rect 8941 9605 8953 9608
rect 8987 9605 8999 9639
rect 9048 9636 9076 9676
rect 9214 9664 9220 9716
rect 9272 9704 9278 9716
rect 10502 9704 10508 9716
rect 9272 9676 10508 9704
rect 9272 9664 9278 9676
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 9122 9636 9128 9648
rect 9048 9608 9128 9636
rect 8941 9599 8999 9605
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 10318 9636 10324 9648
rect 9508 9608 10324 9636
rect 8110 9528 8116 9580
rect 8168 9568 8174 9580
rect 9508 9568 9536 9608
rect 10318 9596 10324 9608
rect 10376 9596 10382 9648
rect 8168 9540 9536 9568
rect 9585 9571 9643 9577
rect 8168 9528 8174 9540
rect 9585 9537 9597 9571
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 9398 9500 9404 9512
rect 7791 9472 9404 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 6052 9404 6408 9432
rect 6052 9392 6058 9404
rect 7834 9392 7840 9444
rect 7892 9432 7898 9444
rect 7892 9404 8340 9432
rect 7892 9392 7898 9404
rect 4120 9336 5212 9364
rect 4120 9324 4126 9336
rect 5810 9324 5816 9376
rect 5868 9324 5874 9376
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9364 6423 9367
rect 6822 9364 6828 9376
rect 6411 9336 6828 9364
rect 6411 9333 6423 9336
rect 6365 9327 6423 9333
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 8018 9324 8024 9376
rect 8076 9324 8082 9376
rect 8202 9324 8208 9376
rect 8260 9324 8266 9376
rect 8312 9364 8340 9404
rect 8570 9392 8576 9444
rect 8628 9392 8634 9444
rect 8757 9435 8815 9441
rect 8757 9401 8769 9435
rect 8803 9401 8815 9435
rect 8757 9395 8815 9401
rect 8772 9364 8800 9395
rect 9214 9392 9220 9444
rect 9272 9432 9278 9444
rect 9309 9435 9367 9441
rect 9309 9432 9321 9435
rect 9272 9404 9321 9432
rect 9272 9392 9278 9404
rect 9309 9401 9321 9404
rect 9355 9401 9367 9435
rect 9309 9395 9367 9401
rect 9493 9435 9551 9441
rect 9493 9401 9505 9435
rect 9539 9401 9551 9435
rect 9600 9432 9628 9531
rect 9766 9528 9772 9580
rect 9824 9528 9830 9580
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9568 10011 9571
rect 10042 9568 10048 9580
rect 9999 9540 10048 9568
rect 9999 9537 10011 9540
rect 9953 9531 10011 9537
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 10244 9500 10272 9531
rect 9968 9472 10272 9500
rect 9600 9404 9812 9432
rect 9493 9395 9551 9401
rect 8312 9336 8800 9364
rect 8941 9367 8999 9373
rect 8941 9333 8953 9367
rect 8987 9364 8999 9367
rect 9122 9364 9128 9376
rect 8987 9336 9128 9364
rect 8987 9333 8999 9336
rect 8941 9327 8999 9333
rect 9122 9324 9128 9336
rect 9180 9364 9186 9376
rect 9508 9364 9536 9395
rect 9784 9376 9812 9404
rect 9674 9364 9680 9376
rect 9180 9336 9680 9364
rect 9180 9324 9186 9336
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 9766 9324 9772 9376
rect 9824 9324 9830 9376
rect 9858 9324 9864 9376
rect 9916 9364 9922 9376
rect 9968 9364 9996 9472
rect 9916 9336 9996 9364
rect 9916 9324 9922 9336
rect 10134 9324 10140 9376
rect 10192 9324 10198 9376
rect 10410 9324 10416 9376
rect 10468 9324 10474 9376
rect 1104 9274 10764 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 10764 9274
rect 1104 9200 10764 9222
rect 3053 9163 3111 9169
rect 3053 9129 3065 9163
rect 3099 9160 3111 9163
rect 3099 9132 6960 9160
rect 3099 9129 3111 9132
rect 3053 9123 3111 9129
rect 1210 9052 1216 9104
rect 1268 9092 1274 9104
rect 4798 9092 4804 9104
rect 1268 9064 4804 9092
rect 1268 9052 1274 9064
rect 4798 9052 4804 9064
rect 4856 9052 4862 9104
rect 6932 9092 6960 9132
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 7837 9163 7895 9169
rect 7837 9160 7849 9163
rect 7708 9132 7849 9160
rect 7708 9120 7714 9132
rect 7837 9129 7849 9132
rect 7883 9129 7895 9163
rect 7837 9123 7895 9129
rect 8294 9120 8300 9172
rect 8352 9120 8358 9172
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 9214 9160 9220 9172
rect 8444 9132 9220 9160
rect 8444 9120 8450 9132
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 10042 9120 10048 9172
rect 10100 9120 10106 9172
rect 8312 9092 8340 9120
rect 6932 9064 8340 9092
rect 2866 8984 2872 9036
rect 2924 9024 2930 9036
rect 2924 8996 3188 9024
rect 2924 8984 2930 8996
rect 2314 8848 2320 8900
rect 2372 8888 2378 8900
rect 2685 8891 2743 8897
rect 2685 8888 2697 8891
rect 2372 8860 2697 8888
rect 2372 8848 2378 8860
rect 2685 8857 2697 8860
rect 2731 8857 2743 8891
rect 2685 8851 2743 8857
rect 2869 8891 2927 8897
rect 2869 8857 2881 8891
rect 2915 8857 2927 8891
rect 3160 8888 3188 8996
rect 3234 8984 3240 9036
rect 3292 9024 3298 9036
rect 3418 9024 3424 9036
rect 3292 8996 3424 9024
rect 3292 8984 3298 8996
rect 3418 8984 3424 8996
rect 3476 9024 3482 9036
rect 5810 9024 5816 9036
rect 3476 8996 5816 9024
rect 3476 8984 3482 8996
rect 4172 8965 4200 8996
rect 5810 8984 5816 8996
rect 5868 8984 5874 9036
rect 7282 8984 7288 9036
rect 7340 9024 7346 9036
rect 9769 9027 9827 9033
rect 9769 9024 9781 9027
rect 7340 8996 8248 9024
rect 7340 8984 7346 8996
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8956 4491 8959
rect 5902 8956 5908 8968
rect 4479 8928 5908 8956
rect 4479 8925 4491 8928
rect 4433 8919 4491 8925
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8956 6055 8959
rect 6638 8956 6644 8968
rect 6043 8928 6644 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 7745 8959 7803 8965
rect 6788 8928 7696 8956
rect 6788 8916 6794 8928
rect 3418 8888 3424 8900
rect 3160 8860 3424 8888
rect 2869 8851 2927 8857
rect 2884 8820 2912 8851
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 4249 8891 4307 8897
rect 4249 8857 4261 8891
rect 4295 8888 4307 8891
rect 4890 8888 4896 8900
rect 4295 8860 4896 8888
rect 4295 8857 4307 8860
rect 4249 8851 4307 8857
rect 4890 8848 4896 8860
rect 4948 8848 4954 8900
rect 5074 8848 5080 8900
rect 5132 8888 5138 8900
rect 5132 8860 5488 8888
rect 5132 8848 5138 8860
rect 4338 8820 4344 8832
rect 2884 8792 4344 8820
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 4617 8823 4675 8829
rect 4617 8789 4629 8823
rect 4663 8820 4675 8823
rect 5350 8820 5356 8832
rect 4663 8792 5356 8820
rect 4663 8789 4675 8792
rect 4617 8783 4675 8789
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 5460 8820 5488 8860
rect 5534 8848 5540 8900
rect 5592 8888 5598 8900
rect 6242 8891 6300 8897
rect 6242 8888 6254 8891
rect 5592 8860 6254 8888
rect 5592 8848 5598 8860
rect 6242 8857 6254 8860
rect 6288 8857 6300 8891
rect 6242 8851 6300 8857
rect 6380 8860 7604 8888
rect 6380 8820 6408 8860
rect 5460 8792 6408 8820
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7576 8829 7604 8860
rect 7377 8823 7435 8829
rect 7377 8820 7389 8823
rect 6972 8792 7389 8820
rect 6972 8780 6978 8792
rect 7377 8789 7389 8792
rect 7423 8789 7435 8823
rect 7377 8783 7435 8789
rect 7561 8823 7619 8829
rect 7561 8789 7573 8823
rect 7607 8789 7619 8823
rect 7668 8820 7696 8928
rect 7745 8925 7757 8959
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 7760 8888 7788 8919
rect 8018 8916 8024 8968
rect 8076 8916 8082 8968
rect 8220 8965 8248 8996
rect 8312 8996 9781 9024
rect 8312 8968 8340 8996
rect 9769 8993 9781 8996
rect 9815 8993 9827 9027
rect 9769 8987 9827 8993
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8294 8916 8300 8968
rect 8352 8916 8358 8968
rect 9214 8916 9220 8968
rect 9272 8956 9278 8968
rect 9582 8956 9588 8968
rect 9272 8928 9588 8956
rect 9272 8916 9278 8928
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 10008 8928 10272 8956
rect 10008 8916 10014 8928
rect 10244 8900 10272 8928
rect 8110 8888 8116 8900
rect 7760 8860 8116 8888
rect 8110 8848 8116 8860
rect 8168 8848 8174 8900
rect 9401 8891 9459 8897
rect 9401 8888 9413 8891
rect 8220 8860 9413 8888
rect 8220 8820 8248 8860
rect 9401 8857 9413 8860
rect 9447 8857 9459 8891
rect 9401 8851 9459 8857
rect 10226 8848 10232 8900
rect 10284 8848 10290 8900
rect 7668 8792 8248 8820
rect 7561 8783 7619 8789
rect 8386 8780 8392 8832
rect 8444 8780 8450 8832
rect 9490 8780 9496 8832
rect 9548 8780 9554 8832
rect 9858 8780 9864 8832
rect 9916 8780 9922 8832
rect 10029 8823 10087 8829
rect 10029 8789 10041 8823
rect 10075 8820 10087 8823
rect 10134 8820 10140 8832
rect 10075 8792 10140 8820
rect 10075 8789 10087 8792
rect 10029 8783 10087 8789
rect 10134 8780 10140 8792
rect 10192 8780 10198 8832
rect 1104 8730 10764 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 7610 8730
rect 7662 8678 7674 8730
rect 7726 8678 7738 8730
rect 7790 8678 7802 8730
rect 7854 8678 7866 8730
rect 7918 8678 10764 8730
rect 1104 8656 10764 8678
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8616 2835 8619
rect 3418 8616 3424 8628
rect 2823 8588 3424 8616
rect 2823 8585 2835 8588
rect 2777 8579 2835 8585
rect 3418 8576 3424 8588
rect 3476 8616 3482 8628
rect 3970 8616 3976 8628
rect 3476 8588 3976 8616
rect 3476 8576 3482 8588
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4246 8576 4252 8628
rect 4304 8616 4310 8628
rect 4817 8619 4875 8625
rect 4817 8616 4829 8619
rect 4304 8588 4829 8616
rect 4304 8576 4310 8588
rect 4817 8585 4829 8588
rect 4863 8585 4875 8619
rect 4817 8579 4875 8585
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 8389 8619 8447 8625
rect 8389 8616 8401 8619
rect 5960 8588 8401 8616
rect 5960 8576 5966 8588
rect 8389 8585 8401 8588
rect 8435 8616 8447 8619
rect 8478 8616 8484 8628
rect 8435 8588 8484 8616
rect 8435 8585 8447 8588
rect 8389 8579 8447 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 10019 8619 10077 8625
rect 10019 8616 10031 8619
rect 8996 8588 10031 8616
rect 8996 8576 9002 8588
rect 10019 8585 10031 8588
rect 10065 8585 10077 8619
rect 10019 8579 10077 8585
rect 4617 8551 4675 8557
rect 1412 8520 4108 8548
rect 1412 8489 1440 8520
rect 1397 8483 1455 8489
rect 1397 8449 1409 8483
rect 1443 8449 1455 8483
rect 1664 8483 1722 8489
rect 1664 8480 1676 8483
rect 1397 8443 1455 8449
rect 1504 8452 1676 8480
rect 1118 8372 1124 8424
rect 1176 8412 1182 8424
rect 1504 8412 1532 8452
rect 1664 8449 1676 8452
rect 1710 8449 1722 8483
rect 1664 8443 1722 8449
rect 4080 8424 4108 8520
rect 4617 8517 4629 8551
rect 4663 8548 4675 8551
rect 4706 8548 4712 8560
rect 4663 8520 4712 8548
rect 4663 8517 4675 8520
rect 4617 8511 4675 8517
rect 4706 8508 4712 8520
rect 4764 8548 4770 8560
rect 10229 8551 10287 8557
rect 4764 8520 9168 8548
rect 4764 8508 4770 8520
rect 9140 8492 9168 8520
rect 10229 8517 10241 8551
rect 10275 8548 10287 8551
rect 10275 8520 10456 8548
rect 10275 8517 10287 8520
rect 10229 8511 10287 8517
rect 5166 8440 5172 8492
rect 5224 8480 5230 8492
rect 5721 8483 5779 8489
rect 5721 8480 5733 8483
rect 5224 8452 5733 8480
rect 5224 8440 5230 8452
rect 5721 8449 5733 8452
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 5994 8440 6000 8492
rect 6052 8440 6058 8492
rect 9122 8440 9128 8492
rect 9180 8440 9186 8492
rect 9513 8483 9571 8489
rect 9513 8449 9525 8483
rect 9559 8480 9571 8483
rect 9674 8480 9680 8492
rect 9559 8452 9680 8480
rect 9559 8449 9571 8452
rect 9513 8443 9571 8449
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 1176 8384 1532 8412
rect 1176 8372 1182 8384
rect 3142 8372 3148 8424
rect 3200 8372 3206 8424
rect 4062 8372 4068 8424
rect 4120 8372 4126 8424
rect 4338 8372 4344 8424
rect 4396 8412 4402 8424
rect 6012 8412 6040 8440
rect 4396 8384 6040 8412
rect 9769 8415 9827 8421
rect 4396 8372 4402 8384
rect 9769 8381 9781 8415
rect 9815 8381 9827 8415
rect 9769 8375 9827 8381
rect 3160 8344 3188 8372
rect 3160 8316 4108 8344
rect 4080 8276 4108 8316
rect 4154 8304 4160 8356
rect 4212 8344 4218 8356
rect 4522 8344 4528 8356
rect 4212 8316 4528 8344
rect 4212 8304 4218 8316
rect 4522 8304 4528 8316
rect 4580 8304 4586 8356
rect 6914 8344 6920 8356
rect 4632 8316 5948 8344
rect 4632 8276 4660 8316
rect 4080 8248 4660 8276
rect 4798 8236 4804 8288
rect 4856 8236 4862 8288
rect 4985 8279 5043 8285
rect 4985 8245 4997 8279
rect 5031 8276 5043 8279
rect 5442 8276 5448 8288
rect 5031 8248 5448 8276
rect 5031 8245 5043 8248
rect 4985 8239 5043 8245
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 5534 8236 5540 8288
rect 5592 8236 5598 8288
rect 5920 8276 5948 8316
rect 6104 8316 6920 8344
rect 6104 8276 6132 8316
rect 6914 8304 6920 8316
rect 6972 8344 6978 8356
rect 8294 8344 8300 8356
rect 6972 8316 8300 8344
rect 6972 8304 6978 8316
rect 8294 8304 8300 8316
rect 8352 8304 8358 8356
rect 5920 8248 6132 8276
rect 9398 8236 9404 8288
rect 9456 8276 9462 8288
rect 9784 8276 9812 8375
rect 9858 8304 9864 8356
rect 9916 8304 9922 8356
rect 10428 8288 10456 8520
rect 9456 8248 9812 8276
rect 9456 8236 9462 8248
rect 10042 8236 10048 8288
rect 10100 8236 10106 8288
rect 10410 8236 10416 8288
rect 10468 8236 10474 8288
rect 1104 8186 10764 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 10764 8186
rect 1104 8112 10764 8134
rect 4890 8072 4896 8084
rect 3896 8044 4896 8072
rect 3896 8013 3924 8044
rect 4890 8032 4896 8044
rect 4948 8032 4954 8084
rect 5258 8032 5264 8084
rect 5316 8072 5322 8084
rect 5537 8075 5595 8081
rect 5537 8072 5549 8075
rect 5316 8044 5549 8072
rect 5316 8032 5322 8044
rect 5537 8041 5549 8044
rect 5583 8072 5595 8075
rect 8754 8072 8760 8084
rect 5583 8044 8760 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 8938 8072 8944 8084
rect 8864 8044 8944 8072
rect 3881 8007 3939 8013
rect 3881 8004 3893 8007
rect 1320 7976 3893 8004
rect 1320 7948 1348 7976
rect 3881 7973 3893 7976
rect 3927 7973 3939 8007
rect 3881 7967 3939 7973
rect 1302 7896 1308 7948
rect 1360 7896 1366 7948
rect 7282 7936 7288 7948
rect 5184 7908 7288 7936
rect 5005 7871 5063 7877
rect 5005 7837 5017 7871
rect 5051 7868 5063 7871
rect 5184 7868 5212 7908
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 8294 7936 8300 7948
rect 7383 7908 8300 7936
rect 5051 7840 5212 7868
rect 5051 7837 5063 7840
rect 5005 7831 5063 7837
rect 5258 7828 5264 7880
rect 5316 7828 5322 7880
rect 5350 7828 5356 7880
rect 5408 7828 5414 7880
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7868 5963 7871
rect 6178 7868 6184 7880
rect 5951 7840 6184 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 6178 7828 6184 7840
rect 6236 7868 6242 7880
rect 6546 7868 6552 7880
rect 6236 7840 6552 7868
rect 6236 7828 6242 7840
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 7383 7868 7411 7908
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 8864 7936 8892 8044
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 8812 7908 8892 7936
rect 8812 7896 8818 7908
rect 8938 7896 8944 7948
rect 8996 7936 9002 7948
rect 8996 7908 9444 7936
rect 8996 7896 9002 7908
rect 6788 7840 7411 7868
rect 6788 7828 6794 7840
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 9416 7877 9444 7908
rect 9401 7871 9459 7877
rect 8720 7864 8800 7868
rect 8720 7844 9076 7864
rect 9125 7849 9183 7855
rect 9125 7844 9137 7849
rect 8720 7840 9137 7844
rect 8720 7828 8726 7840
rect 8772 7836 9137 7840
rect 4890 7800 4896 7812
rect 2976 7772 4896 7800
rect 2976 7744 3004 7772
rect 4890 7760 4896 7772
rect 4948 7760 4954 7812
rect 5368 7800 5396 7828
rect 9048 7816 9137 7836
rect 9125 7815 9137 7816
rect 9171 7815 9183 7849
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7868 10287 7871
rect 10410 7868 10416 7880
rect 10275 7840 10416 7868
rect 10275 7837 10287 7840
rect 10229 7831 10287 7837
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 5537 7803 5595 7809
rect 5537 7800 5549 7803
rect 5368 7772 5549 7800
rect 5537 7769 5549 7772
rect 5583 7769 5595 7803
rect 5537 7763 5595 7769
rect 6086 7760 6092 7812
rect 6144 7800 6150 7812
rect 6638 7800 6644 7812
rect 6144 7772 6644 7800
rect 6144 7760 6150 7772
rect 6638 7760 6644 7772
rect 6696 7760 6702 7812
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 8294 7800 8300 7812
rect 6972 7772 8300 7800
rect 6972 7760 6978 7772
rect 8294 7760 8300 7772
rect 8352 7760 8358 7812
rect 9125 7809 9183 7815
rect 9585 7803 9643 7809
rect 9585 7769 9597 7803
rect 9631 7800 9643 7803
rect 10594 7800 10600 7812
rect 9631 7772 10600 7800
rect 9631 7769 9643 7772
rect 9585 7763 9643 7769
rect 10594 7760 10600 7772
rect 10652 7760 10658 7812
rect 2958 7692 2964 7744
rect 3016 7692 3022 7744
rect 3418 7692 3424 7744
rect 3476 7732 3482 7744
rect 3694 7732 3700 7744
rect 3476 7704 3700 7732
rect 3476 7692 3482 7704
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 5350 7692 5356 7744
rect 5408 7692 5414 7744
rect 5626 7692 5632 7744
rect 5684 7732 5690 7744
rect 8754 7732 8760 7744
rect 5684 7704 8760 7732
rect 5684 7692 5690 7704
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 9214 7692 9220 7744
rect 9272 7692 9278 7744
rect 10410 7692 10416 7744
rect 10468 7692 10474 7744
rect 1104 7642 10764 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 10764 7642
rect 1104 7568 10764 7590
rect 2498 7488 2504 7540
rect 2556 7528 2562 7540
rect 2685 7531 2743 7537
rect 2685 7528 2697 7531
rect 2556 7500 2697 7528
rect 2556 7488 2562 7500
rect 2685 7497 2697 7500
rect 2731 7528 2743 7531
rect 3694 7528 3700 7540
rect 2731 7500 3700 7528
rect 2731 7497 2743 7500
rect 2685 7491 2743 7497
rect 3694 7488 3700 7500
rect 3752 7488 3758 7540
rect 3970 7488 3976 7540
rect 4028 7488 4034 7540
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 6549 7531 6607 7537
rect 5500 7500 6408 7528
rect 5500 7488 5506 7500
rect 3050 7460 3056 7472
rect 2746 7432 3056 7460
rect 2746 7404 2774 7432
rect 3050 7420 3056 7432
rect 3108 7460 3114 7472
rect 3988 7460 4016 7488
rect 3108 7432 4016 7460
rect 4976 7463 5034 7469
rect 3108 7420 3114 7432
rect 4976 7429 4988 7463
rect 5022 7460 5034 7463
rect 5534 7460 5540 7472
rect 5022 7432 5540 7460
rect 5022 7429 5034 7432
rect 4976 7423 5034 7429
rect 5534 7420 5540 7432
rect 5592 7420 5598 7472
rect 1486 7352 1492 7404
rect 1544 7352 1550 7404
rect 2682 7352 2688 7404
rect 2740 7364 2774 7404
rect 3809 7395 3867 7401
rect 2740 7352 2746 7364
rect 3809 7361 3821 7395
rect 3855 7392 3867 7395
rect 4154 7392 4160 7404
rect 3855 7364 4160 7392
rect 3855 7361 3867 7364
rect 3809 7355 3867 7361
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 6380 7401 6408 7500
rect 6549 7497 6561 7531
rect 6595 7528 6607 7531
rect 7466 7528 7472 7540
rect 6595 7500 7472 7528
rect 6595 7497 6607 7500
rect 6549 7491 6607 7497
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8938 7528 8944 7540
rect 8260 7500 8944 7528
rect 8260 7488 8266 7500
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 9769 7531 9827 7537
rect 9769 7497 9781 7531
rect 9815 7528 9827 7531
rect 10318 7528 10324 7540
rect 9815 7500 10324 7528
rect 9815 7497 9827 7500
rect 9769 7491 9827 7497
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 7374 7420 7380 7472
rect 7432 7460 7438 7472
rect 9953 7463 10011 7469
rect 9953 7460 9965 7463
rect 7432 7432 9965 7460
rect 7432 7420 7438 7432
rect 9953 7429 9965 7432
rect 9999 7429 10011 7463
rect 9953 7423 10011 7429
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7392 4675 7395
rect 6365 7395 6423 7401
rect 4663 7364 5948 7392
rect 4663 7361 4675 7364
rect 4617 7355 4675 7361
rect 4062 7284 4068 7336
rect 4120 7324 4126 7336
rect 4709 7327 4767 7333
rect 4709 7324 4721 7327
rect 4120 7296 4721 7324
rect 4120 7284 4126 7296
rect 4709 7293 4721 7296
rect 4755 7293 4767 7327
rect 4709 7287 4767 7293
rect 5920 7200 5948 7364
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 6880 7364 7941 7392
rect 6880 7352 6886 7364
rect 7929 7361 7941 7364
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 10594 7392 10600 7404
rect 8352 7364 10600 7392
rect 8352 7352 8358 7364
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 5994 7284 6000 7336
rect 6052 7324 6058 7336
rect 9490 7324 9496 7336
rect 6052 7296 9496 7324
rect 6052 7284 6058 7296
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 6089 7259 6147 7265
rect 6089 7225 6101 7259
rect 6135 7256 6147 7259
rect 6638 7256 6644 7268
rect 6135 7228 6644 7256
rect 6135 7225 6147 7228
rect 6089 7219 6147 7225
rect 6638 7216 6644 7228
rect 6696 7256 6702 7268
rect 8938 7256 8944 7268
rect 6696 7228 8944 7256
rect 6696 7216 6702 7228
rect 8938 7216 8944 7228
rect 8996 7216 9002 7268
rect 9306 7216 9312 7268
rect 9364 7256 9370 7268
rect 9364 7228 9996 7256
rect 9364 7216 9370 7228
rect 750 7148 756 7200
rect 808 7188 814 7200
rect 1581 7191 1639 7197
rect 1581 7188 1593 7191
rect 808 7160 1593 7188
rect 808 7148 814 7160
rect 1581 7157 1593 7160
rect 1627 7157 1639 7191
rect 1581 7151 1639 7157
rect 4525 7191 4583 7197
rect 4525 7157 4537 7191
rect 4571 7188 4583 7191
rect 4614 7188 4620 7200
rect 4571 7160 4620 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 5902 7148 5908 7200
rect 5960 7188 5966 7200
rect 7558 7188 7564 7200
rect 5960 7160 7564 7188
rect 5960 7148 5966 7160
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 8754 7148 8760 7200
rect 8812 7188 8818 7200
rect 9217 7191 9275 7197
rect 9217 7188 9229 7191
rect 8812 7160 9229 7188
rect 8812 7148 8818 7160
rect 9217 7157 9229 7160
rect 9263 7188 9275 7191
rect 9398 7188 9404 7200
rect 9263 7160 9404 7188
rect 9263 7157 9275 7160
rect 9217 7151 9275 7157
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 9968 7197 9996 7228
rect 10318 7216 10324 7268
rect 10376 7216 10382 7268
rect 9953 7191 10011 7197
rect 9953 7157 9965 7191
rect 9999 7157 10011 7191
rect 9953 7151 10011 7157
rect 1104 7098 10764 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 10764 7098
rect 1104 7024 10764 7046
rect 2682 6984 2688 6996
rect 1780 6956 2688 6984
rect 1780 6789 1808 6956
rect 2682 6944 2688 6956
rect 2740 6984 2746 6996
rect 3421 6987 3479 6993
rect 3421 6984 3433 6987
rect 2740 6956 3433 6984
rect 2740 6944 2746 6956
rect 3421 6953 3433 6956
rect 3467 6953 3479 6987
rect 3421 6947 3479 6953
rect 3786 6944 3792 6996
rect 3844 6944 3850 6996
rect 4264 6956 5212 6984
rect 2222 6876 2228 6928
rect 2280 6916 2286 6928
rect 4264 6916 4292 6956
rect 2280 6888 4292 6916
rect 5184 6916 5212 6956
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 6822 6984 6828 6996
rect 5592 6956 6828 6984
rect 5592 6944 5598 6956
rect 6822 6944 6828 6956
rect 6880 6984 6886 6996
rect 6917 6987 6975 6993
rect 6917 6984 6929 6987
rect 6880 6956 6929 6984
rect 6880 6944 6886 6956
rect 6917 6953 6929 6956
rect 6963 6953 6975 6987
rect 6917 6947 6975 6953
rect 7374 6944 7380 6996
rect 7432 6984 7438 6996
rect 8662 6984 8668 6996
rect 7432 6956 8668 6984
rect 7432 6944 7438 6956
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 10042 6944 10048 6996
rect 10100 6944 10106 6996
rect 10060 6916 10088 6944
rect 5184 6888 10088 6916
rect 2280 6876 2286 6888
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6848 2375 6851
rect 2498 6848 2504 6860
rect 2363 6820 2504 6848
rect 2363 6817 2375 6820
rect 2317 6811 2375 6817
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 2792 6820 3188 6848
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6749 1823 6783
rect 1765 6743 1823 6749
rect 1946 6740 1952 6792
rect 2004 6740 2010 6792
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6749 2099 6783
rect 2041 6743 2099 6749
rect 2133 6783 2191 6789
rect 2133 6749 2145 6783
rect 2179 6749 2191 6783
rect 2133 6743 2191 6749
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6780 2651 6783
rect 2682 6780 2688 6792
rect 2639 6752 2688 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 1946 6644 1952 6656
rect 1627 6616 1952 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 1946 6604 1952 6616
rect 2004 6604 2010 6656
rect 2056 6644 2084 6743
rect 2148 6712 2176 6743
rect 2682 6740 2688 6752
rect 2740 6740 2746 6792
rect 2792 6712 2820 6820
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 3160 6780 3188 6820
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 3878 6848 3884 6860
rect 3292 6820 3884 6848
rect 3292 6808 3298 6820
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 5902 6848 5908 6860
rect 5092 6820 5908 6848
rect 3326 6780 3332 6792
rect 3160 6752 3332 6780
rect 2869 6743 2927 6749
rect 2148 6684 2820 6712
rect 2130 6644 2136 6656
rect 2056 6616 2136 6644
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 2314 6604 2320 6656
rect 2372 6604 2378 6656
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 2590 6644 2596 6656
rect 2455 6616 2596 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 2590 6604 2596 6616
rect 2648 6604 2654 6656
rect 2774 6604 2780 6656
rect 2832 6604 2838 6656
rect 2884 6644 2912 6743
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 5092 6780 5120 6820
rect 5902 6808 5908 6820
rect 5960 6848 5966 6860
rect 6362 6848 6368 6860
rect 5960 6820 6368 6848
rect 5960 6808 5966 6820
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 6638 6808 6644 6860
rect 6696 6848 6702 6860
rect 7374 6848 7380 6860
rect 6696 6820 7380 6848
rect 6696 6808 6702 6820
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 4816 6752 5120 6780
rect 5169 6783 5227 6789
rect 3234 6672 3240 6724
rect 3292 6672 3298 6724
rect 4816 6712 4844 6752
rect 5169 6749 5181 6783
rect 5215 6780 5227 6783
rect 5258 6780 5264 6792
rect 5215 6752 5264 6780
rect 5215 6749 5227 6752
rect 5169 6743 5227 6749
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 6086 6780 6092 6792
rect 5776 6752 6092 6780
rect 5776 6740 5782 6752
rect 6086 6740 6092 6752
rect 6144 6780 6150 6792
rect 8202 6780 8208 6792
rect 6144 6752 8208 6780
rect 6144 6740 6150 6752
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8294 6740 8300 6792
rect 8352 6780 8358 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 8352 6752 8401 6780
rect 8352 6740 8358 6752
rect 8389 6749 8401 6752
rect 8435 6749 8447 6783
rect 9306 6780 9312 6792
rect 8389 6743 8447 6749
rect 8496 6752 9312 6780
rect 3344 6684 4844 6712
rect 4924 6715 4982 6721
rect 3344 6644 3372 6684
rect 4924 6681 4936 6715
rect 4970 6712 4982 6715
rect 4970 6684 5396 6712
rect 4970 6681 4982 6684
rect 4924 6675 4982 6681
rect 2884 6616 3372 6644
rect 3418 6604 3424 6656
rect 3476 6653 3482 6656
rect 3476 6647 3495 6653
rect 3483 6613 3495 6647
rect 3476 6607 3495 6613
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 3694 6644 3700 6656
rect 3651 6616 3700 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 3476 6604 3482 6607
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 5368 6644 5396 6684
rect 5442 6672 5448 6724
rect 5500 6712 5506 6724
rect 5629 6715 5687 6721
rect 5629 6712 5641 6715
rect 5500 6684 5641 6712
rect 5500 6672 5506 6684
rect 5629 6681 5641 6684
rect 5675 6681 5687 6715
rect 5629 6675 5687 6681
rect 6546 6672 6552 6724
rect 6604 6712 6610 6724
rect 8496 6712 8524 6752
rect 9306 6740 9312 6752
rect 9364 6780 9370 6792
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 9364 6752 9505 6780
rect 9364 6740 9370 6752
rect 9493 6749 9505 6752
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 6604 6684 8524 6712
rect 6604 6672 6610 6684
rect 8938 6672 8944 6724
rect 8996 6712 9002 6724
rect 9692 6712 9720 6743
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10134 6712 10140 6724
rect 8996 6684 10140 6712
rect 8996 6672 9002 6684
rect 10134 6672 10140 6684
rect 10192 6672 10198 6724
rect 8205 6647 8263 6653
rect 8205 6644 8217 6647
rect 5368 6616 8217 6644
rect 8205 6613 8217 6616
rect 8251 6613 8263 6647
rect 8205 6607 8263 6613
rect 9582 6604 9588 6656
rect 9640 6604 9646 6656
rect 10410 6604 10416 6656
rect 10468 6604 10474 6656
rect 1104 6554 10764 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 10764 6554
rect 1104 6480 10764 6502
rect 1486 6400 1492 6452
rect 1544 6400 1550 6452
rect 1673 6443 1731 6449
rect 1673 6409 1685 6443
rect 1719 6440 1731 6443
rect 1854 6440 1860 6452
rect 1719 6412 1860 6440
rect 1719 6409 1731 6412
rect 1673 6403 1731 6409
rect 1854 6400 1860 6412
rect 1912 6400 1918 6452
rect 1949 6443 2007 6449
rect 1949 6409 1961 6443
rect 1995 6440 2007 6443
rect 2222 6440 2228 6452
rect 1995 6412 2228 6440
rect 1995 6409 2007 6412
rect 1949 6403 2007 6409
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 2700 6412 3188 6440
rect 1504 6372 1532 6400
rect 2700 6384 2728 6412
rect 1504 6344 1808 6372
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 1780 6313 1808 6344
rect 2682 6332 2688 6384
rect 2740 6332 2746 6384
rect 2866 6332 2872 6384
rect 2924 6381 2930 6384
rect 2924 6375 2959 6381
rect 2947 6341 2959 6375
rect 2924 6335 2959 6341
rect 2924 6332 2930 6335
rect 3160 6313 3188 6412
rect 3252 6412 4660 6440
rect 1489 6307 1547 6313
rect 1489 6304 1501 6307
rect 1360 6276 1501 6304
rect 1360 6264 1366 6276
rect 1489 6273 1501 6276
rect 1535 6273 1547 6307
rect 1489 6267 1547 6273
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6273 3203 6307
rect 3145 6267 3203 6273
rect 1964 6236 1992 6267
rect 3252 6236 3280 6412
rect 4338 6372 4344 6384
rect 3344 6344 4344 6372
rect 3344 6313 3372 6344
rect 4338 6332 4344 6344
rect 4396 6332 4402 6384
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6273 3387 6307
rect 3329 6267 3387 6273
rect 3418 6264 3424 6316
rect 3476 6264 3482 6316
rect 3510 6264 3516 6316
rect 3568 6264 3574 6316
rect 3697 6307 3755 6313
rect 3697 6273 3709 6307
rect 3743 6304 3755 6307
rect 4632 6304 4660 6412
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 5684 6412 5856 6440
rect 5684 6400 5690 6412
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 5721 6375 5779 6381
rect 5721 6372 5733 6375
rect 5592 6344 5733 6372
rect 5592 6332 5598 6344
rect 5721 6341 5733 6344
rect 5767 6341 5779 6375
rect 5721 6335 5779 6341
rect 5828 6304 5856 6412
rect 6012 6412 6316 6440
rect 6012 6381 6040 6412
rect 5997 6375 6055 6381
rect 5997 6341 6009 6375
rect 6043 6341 6055 6375
rect 5997 6335 6055 6341
rect 6086 6332 6092 6384
rect 6144 6372 6150 6384
rect 6181 6375 6239 6381
rect 6181 6372 6193 6375
rect 6144 6344 6193 6372
rect 6144 6332 6150 6344
rect 6181 6341 6193 6344
rect 6227 6341 6239 6375
rect 6288 6372 6316 6412
rect 6454 6400 6460 6452
rect 6512 6400 6518 6452
rect 6638 6440 6644 6452
rect 6564 6412 6644 6440
rect 6564 6372 6592 6412
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 7926 6440 7932 6452
rect 6748 6412 7932 6440
rect 6748 6384 6776 6412
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 8481 6443 8539 6449
rect 8481 6440 8493 6443
rect 8260 6412 8493 6440
rect 8260 6400 8266 6412
rect 8481 6409 8493 6412
rect 8527 6409 8539 6443
rect 8481 6403 8539 6409
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 8849 6443 8907 6449
rect 8849 6440 8861 6443
rect 8720 6412 8861 6440
rect 8720 6400 8726 6412
rect 8849 6409 8861 6412
rect 8895 6409 8907 6443
rect 8849 6403 8907 6409
rect 8938 6400 8944 6452
rect 8996 6400 9002 6452
rect 9122 6400 9128 6452
rect 9180 6440 9186 6452
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 9180 6412 10057 6440
rect 9180 6400 9186 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10318 6440 10324 6452
rect 10045 6403 10103 6409
rect 10152 6412 10324 6440
rect 6730 6372 6736 6384
rect 6288 6344 6592 6372
rect 6656 6344 6736 6372
rect 6181 6335 6239 6341
rect 6656 6313 6684 6344
rect 6730 6332 6736 6344
rect 6788 6332 6794 6384
rect 6914 6332 6920 6384
rect 6972 6332 6978 6384
rect 7368 6375 7426 6381
rect 7368 6341 7380 6375
rect 7414 6372 7426 6375
rect 7650 6372 7656 6384
rect 7414 6344 7656 6372
rect 7414 6341 7426 6344
rect 7368 6335 7426 6341
rect 7650 6332 7656 6344
rect 7708 6332 7714 6384
rect 7742 6332 7748 6384
rect 7800 6372 7806 6384
rect 8573 6375 8631 6381
rect 8573 6372 8585 6375
rect 7800 6344 8585 6372
rect 7800 6332 7806 6344
rect 8573 6341 8585 6344
rect 8619 6372 8631 6375
rect 8619 6344 8892 6372
rect 8619 6341 8631 6344
rect 8573 6335 8631 6341
rect 5905 6307 5963 6313
rect 5905 6306 5917 6307
rect 5904 6304 5917 6306
rect 3743 6276 4108 6304
rect 4632 6276 5917 6304
rect 3743 6273 3755 6276
rect 3697 6267 3755 6273
rect 1504 6208 3280 6236
rect 1504 6180 1532 6208
rect 3786 6196 3792 6248
rect 3844 6236 3850 6248
rect 3970 6236 3976 6248
rect 3844 6208 3976 6236
rect 3844 6196 3850 6208
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 4080 6236 4108 6276
rect 5905 6273 5917 6276
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6273 6699 6307
rect 6932 6304 6960 6332
rect 8757 6307 8815 6313
rect 8757 6304 8769 6307
rect 6932 6302 7308 6304
rect 7484 6302 8769 6304
rect 6932 6276 8769 6302
rect 7280 6274 7512 6276
rect 6641 6267 6699 6273
rect 8757 6273 8769 6276
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 4246 6236 4252 6248
rect 4080 6208 4252 6236
rect 4246 6196 4252 6208
rect 4304 6196 4310 6248
rect 6454 6196 6460 6248
rect 6512 6236 6518 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6512 6208 6837 6236
rect 6512 6196 6518 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 7098 6196 7104 6248
rect 7156 6196 7162 6248
rect 8478 6196 8484 6248
rect 8536 6236 8542 6248
rect 8864 6236 8892 6344
rect 9030 6332 9036 6384
rect 9088 6332 9094 6384
rect 9214 6332 9220 6384
rect 9272 6372 9278 6384
rect 9369 6375 9427 6381
rect 9369 6372 9381 6375
rect 9272 6344 9381 6372
rect 9272 6332 9278 6344
rect 9369 6341 9381 6344
rect 9415 6341 9427 6375
rect 9369 6335 9427 6341
rect 9585 6375 9643 6381
rect 9585 6341 9597 6375
rect 9631 6341 9643 6375
rect 9585 6335 9643 6341
rect 9677 6375 9735 6381
rect 9677 6341 9689 6375
rect 9723 6372 9735 6375
rect 9766 6372 9772 6384
rect 9723 6344 9772 6372
rect 9723 6341 9735 6344
rect 9677 6335 9735 6341
rect 9048 6304 9076 6332
rect 9600 6304 9628 6335
rect 9766 6332 9772 6344
rect 9824 6332 9830 6384
rect 9861 6375 9919 6381
rect 9861 6341 9873 6375
rect 9907 6372 9919 6375
rect 10152 6372 10180 6412
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 9907 6344 10180 6372
rect 9907 6341 9919 6344
rect 9861 6335 9919 6341
rect 10226 6332 10232 6384
rect 10284 6332 10290 6384
rect 9048 6276 9628 6304
rect 8536 6208 8892 6236
rect 8536 6196 8542 6208
rect 9398 6196 9404 6248
rect 9456 6236 9462 6248
rect 9456 6208 9674 6236
rect 9456 6196 9462 6208
rect 1486 6128 1492 6180
rect 1544 6128 1550 6180
rect 5905 6171 5963 6177
rect 5905 6168 5917 6171
rect 2884 6140 5917 6168
rect 2222 6060 2228 6112
rect 2280 6100 2286 6112
rect 2406 6100 2412 6112
rect 2280 6072 2412 6100
rect 2280 6060 2286 6072
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 2884 6109 2912 6140
rect 5905 6137 5917 6140
rect 5951 6137 5963 6171
rect 8570 6168 8576 6180
rect 5905 6131 5963 6137
rect 8266 6140 8576 6168
rect 2869 6103 2927 6109
rect 2869 6069 2881 6103
rect 2915 6069 2927 6103
rect 2869 6063 2927 6069
rect 3053 6103 3111 6109
rect 3053 6069 3065 6103
rect 3099 6100 3111 6103
rect 3786 6100 3792 6112
rect 3099 6072 3792 6100
rect 3099 6069 3111 6072
rect 3053 6063 3111 6069
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 3878 6060 3884 6112
rect 3936 6060 3942 6112
rect 4982 6060 4988 6112
rect 5040 6100 5046 6112
rect 5626 6100 5632 6112
rect 5040 6072 5632 6100
rect 5040 6060 5046 6072
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 8266 6100 8294 6140
rect 8570 6128 8576 6140
rect 8628 6168 8634 6180
rect 9646 6168 9674 6208
rect 10244 6168 10272 6332
rect 8628 6140 9260 6168
rect 9646 6140 10272 6168
rect 8628 6128 8634 6140
rect 5776 6072 8294 6100
rect 5776 6060 5782 6072
rect 8938 6060 8944 6112
rect 8996 6100 9002 6112
rect 9232 6109 9260 6140
rect 9125 6103 9183 6109
rect 9125 6100 9137 6103
rect 8996 6072 9137 6100
rect 8996 6060 9002 6072
rect 9125 6069 9137 6072
rect 9171 6069 9183 6103
rect 9125 6063 9183 6069
rect 9217 6103 9275 6109
rect 9217 6069 9229 6103
rect 9263 6069 9275 6103
rect 9217 6063 9275 6069
rect 9398 6060 9404 6112
rect 9456 6060 9462 6112
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 10318 6100 10324 6112
rect 9548 6072 10324 6100
rect 9548 6060 9554 6072
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 1104 6010 10764 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 10764 6010
rect 1104 5936 10764 5958
rect 1486 5856 1492 5908
rect 1544 5856 1550 5908
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 4709 5899 4767 5905
rect 4709 5896 4721 5899
rect 4212 5868 4721 5896
rect 4212 5856 4218 5868
rect 4709 5865 4721 5868
rect 4755 5865 4767 5899
rect 4709 5859 4767 5865
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 5534 5896 5540 5908
rect 4856 5868 5540 5896
rect 4856 5856 4862 5868
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 5626 5856 5632 5908
rect 5684 5896 5690 5908
rect 6089 5899 6147 5905
rect 6089 5896 6101 5899
rect 5684 5868 6101 5896
rect 5684 5856 5690 5868
rect 6089 5865 6101 5868
rect 6135 5865 6147 5899
rect 6089 5859 6147 5865
rect 6196 5868 6592 5896
rect 3694 5828 3700 5840
rect 2884 5800 3700 5828
rect 2884 5769 2912 5800
rect 3694 5788 3700 5800
rect 3752 5828 3758 5840
rect 5258 5828 5264 5840
rect 3752 5800 5264 5828
rect 3752 5788 3758 5800
rect 5258 5788 5264 5800
rect 5316 5788 5322 5840
rect 5718 5828 5724 5840
rect 5368 5800 5724 5828
rect 2869 5763 2927 5769
rect 2869 5729 2881 5763
rect 2915 5729 2927 5763
rect 2869 5723 2927 5729
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4212 5732 5304 5760
rect 4212 5720 4218 5732
rect 2590 5652 2596 5704
rect 2648 5701 2654 5704
rect 2648 5695 2671 5701
rect 2659 5661 2671 5695
rect 2648 5655 2671 5661
rect 2648 5652 2654 5655
rect 4430 5652 4436 5704
rect 4488 5692 4494 5704
rect 5276 5701 5304 5732
rect 5368 5701 5396 5800
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 6196 5828 6224 5868
rect 6120 5800 6224 5828
rect 6273 5831 6331 5837
rect 4893 5695 4951 5701
rect 4893 5692 4905 5695
rect 4488 5664 4905 5692
rect 4488 5652 4494 5664
rect 4893 5661 4905 5664
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5661 5319 5695
rect 5261 5655 5319 5661
rect 5353 5695 5411 5701
rect 5353 5661 5365 5695
rect 5399 5661 5411 5695
rect 5353 5655 5411 5661
rect 5445 5695 5503 5701
rect 5445 5661 5457 5695
rect 5491 5692 5503 5695
rect 5718 5692 5724 5704
rect 5491 5664 5724 5692
rect 5491 5661 5503 5664
rect 5445 5655 5503 5661
rect 3510 5584 3516 5636
rect 3568 5624 3574 5636
rect 3568 5596 4568 5624
rect 3568 5584 3574 5596
rect 2682 5516 2688 5568
rect 2740 5556 2746 5568
rect 4430 5556 4436 5568
rect 2740 5528 4436 5556
rect 2740 5516 2746 5528
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 4540 5556 4568 5596
rect 4706 5584 4712 5636
rect 4764 5624 4770 5636
rect 5092 5624 5120 5655
rect 4764 5596 5120 5624
rect 4764 5584 4770 5596
rect 5460 5556 5488 5655
rect 5718 5652 5724 5664
rect 5776 5652 5782 5704
rect 5905 5627 5963 5633
rect 5905 5593 5917 5627
rect 5951 5624 5963 5627
rect 6120 5624 6148 5800
rect 6273 5797 6285 5831
rect 6319 5797 6331 5831
rect 6564 5828 6592 5868
rect 7374 5856 7380 5908
rect 7432 5856 7438 5908
rect 10042 5896 10048 5908
rect 9324 5868 10048 5896
rect 7098 5828 7104 5840
rect 6564 5800 7104 5828
rect 6273 5791 6331 5797
rect 6178 5720 6184 5772
rect 6236 5720 6242 5772
rect 6288 5760 6316 5791
rect 7098 5788 7104 5800
rect 7156 5788 7162 5840
rect 8938 5788 8944 5840
rect 8996 5828 9002 5840
rect 9324 5828 9352 5868
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 8996 5800 9352 5828
rect 8996 5788 9002 5800
rect 9398 5788 9404 5840
rect 9456 5788 9462 5840
rect 9493 5831 9551 5837
rect 9493 5797 9505 5831
rect 9539 5828 9551 5831
rect 10226 5828 10232 5840
rect 9539 5800 10232 5828
rect 9539 5797 9551 5800
rect 9493 5791 9551 5797
rect 10226 5788 10232 5800
rect 10284 5788 10290 5840
rect 6546 5760 6552 5772
rect 6288 5732 6552 5760
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 9030 5760 9036 5772
rect 6656 5732 7420 5760
rect 6196 5692 6224 5720
rect 6656 5701 6684 5732
rect 6365 5695 6423 5701
rect 6365 5692 6377 5695
rect 6196 5664 6377 5692
rect 6365 5661 6377 5664
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 5951 5596 6148 5624
rect 5951 5593 5963 5596
rect 5905 5587 5963 5593
rect 6270 5584 6276 5636
rect 6328 5624 6334 5636
rect 6656 5624 6684 5655
rect 6914 5652 6920 5704
rect 6972 5652 6978 5704
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 7101 5695 7159 5701
rect 7101 5692 7113 5695
rect 7064 5664 7113 5692
rect 7064 5652 7070 5664
rect 7101 5661 7113 5664
rect 7147 5661 7159 5695
rect 7392 5692 7420 5732
rect 8680 5732 9036 5760
rect 8680 5692 8708 5732
rect 9030 5720 9036 5732
rect 9088 5760 9094 5772
rect 9088 5732 10272 5760
rect 9088 5720 9094 5732
rect 7392 5664 8708 5692
rect 7101 5655 7159 5661
rect 8754 5652 8760 5704
rect 8812 5652 8818 5704
rect 8846 5652 8852 5704
rect 8904 5652 8910 5704
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5692 9183 5695
rect 9214 5692 9220 5704
rect 9171 5664 9220 5692
rect 9171 5661 9183 5664
rect 9125 5655 9183 5661
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5692 9735 5695
rect 9858 5692 9864 5704
rect 9723 5664 9864 5692
rect 9723 5661 9735 5664
rect 9677 5655 9735 5661
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 10244 5701 10272 5732
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5661 10287 5695
rect 10229 5655 10287 5661
rect 6328 5596 6684 5624
rect 6825 5627 6883 5633
rect 6328 5584 6334 5596
rect 6825 5593 6837 5627
rect 6871 5593 6883 5627
rect 6825 5587 6883 5593
rect 4540 5528 5488 5556
rect 5718 5516 5724 5568
rect 5776 5516 5782 5568
rect 5810 5516 5816 5568
rect 5868 5556 5874 5568
rect 6086 5556 6092 5568
rect 6144 5565 6150 5568
rect 6144 5559 6163 5565
rect 5868 5528 6092 5556
rect 5868 5516 5874 5528
rect 6086 5516 6092 5528
rect 6151 5525 6163 5559
rect 6144 5519 6163 5525
rect 6144 5516 6150 5519
rect 6454 5516 6460 5568
rect 6512 5516 6518 5568
rect 6730 5516 6736 5568
rect 6788 5556 6794 5568
rect 6840 5556 6868 5587
rect 7374 5584 7380 5636
rect 7432 5624 7438 5636
rect 7650 5624 7656 5636
rect 7432 5596 7656 5624
rect 7432 5584 7438 5596
rect 7650 5584 7656 5596
rect 7708 5584 7714 5636
rect 7742 5584 7748 5636
rect 7800 5584 7806 5636
rect 8018 5584 8024 5636
rect 8076 5584 8082 5636
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 8490 5627 8548 5633
rect 8490 5624 8502 5627
rect 8444 5596 8502 5624
rect 8444 5584 8450 5596
rect 8490 5593 8502 5596
rect 8536 5593 8548 5627
rect 8772 5624 8800 5652
rect 8490 5587 8548 5593
rect 8680 5596 8800 5624
rect 8864 5624 8892 5652
rect 9401 5627 9459 5633
rect 9401 5624 9413 5627
rect 8864 5596 9413 5624
rect 6788 5528 6868 5556
rect 6788 5516 6794 5528
rect 6914 5516 6920 5568
rect 6972 5516 6978 5568
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 7760 5556 7788 5584
rect 7156 5528 7788 5556
rect 8036 5556 8064 5584
rect 8680 5568 8708 5596
rect 9401 5593 9413 5596
rect 9447 5593 9459 5627
rect 9401 5587 9459 5593
rect 8570 5556 8576 5568
rect 8036 5528 8576 5556
rect 7156 5516 7162 5528
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 8662 5516 8668 5568
rect 8720 5516 8726 5568
rect 9214 5516 9220 5568
rect 9272 5516 9278 5568
rect 9490 5516 9496 5568
rect 9548 5556 9554 5568
rect 9858 5556 9864 5568
rect 9548 5528 9864 5556
rect 9548 5516 9554 5528
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 10410 5516 10416 5568
rect 10468 5516 10474 5568
rect 1104 5466 10764 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 10764 5466
rect 1104 5392 10764 5414
rect 1946 5312 1952 5364
rect 2004 5312 2010 5364
rect 5442 5352 5448 5364
rect 2746 5324 5448 5352
rect 1765 5287 1823 5293
rect 1765 5253 1777 5287
rect 1811 5284 1823 5287
rect 2746 5284 2774 5324
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 5534 5312 5540 5364
rect 5592 5312 5598 5364
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 5721 5355 5779 5361
rect 5721 5352 5733 5355
rect 5684 5324 5733 5352
rect 5684 5312 5690 5324
rect 5721 5321 5733 5324
rect 5767 5321 5779 5355
rect 5721 5315 5779 5321
rect 5889 5355 5947 5361
rect 5889 5321 5901 5355
rect 5935 5352 5947 5355
rect 5994 5352 6000 5364
rect 5935 5324 6000 5352
rect 5935 5321 5947 5324
rect 5889 5315 5947 5321
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 10111 5355 10169 5361
rect 10111 5352 10123 5355
rect 6932 5324 10123 5352
rect 6932 5296 6960 5324
rect 10111 5321 10123 5324
rect 10157 5321 10169 5355
rect 10111 5315 10169 5321
rect 1811 5256 2774 5284
rect 2869 5287 2927 5293
rect 1811 5253 1823 5256
rect 1765 5247 1823 5253
rect 2869 5253 2881 5287
rect 2915 5253 2927 5287
rect 2869 5247 2927 5253
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5216 1455 5219
rect 1486 5216 1492 5228
rect 1443 5188 1492 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 1486 5176 1492 5188
rect 1544 5216 1550 5228
rect 2222 5216 2228 5228
rect 1544 5188 2228 5216
rect 1544 5176 1550 5188
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5185 2743 5219
rect 2884 5216 2912 5247
rect 4062 5244 4068 5296
rect 4120 5284 4126 5296
rect 6089 5287 6147 5293
rect 6089 5284 6101 5287
rect 4120 5256 5396 5284
rect 4120 5244 4126 5256
rect 3142 5216 3148 5228
rect 2884 5188 3148 5216
rect 2685 5179 2743 5185
rect 2700 5148 2728 5179
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 4890 5176 4896 5228
rect 4948 5225 4954 5228
rect 4948 5216 4960 5225
rect 5368 5216 5396 5256
rect 5552 5256 6101 5284
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 4948 5188 4993 5216
rect 5368 5188 5457 5216
rect 4948 5179 4960 5188
rect 4948 5176 4954 5179
rect 2958 5148 2964 5160
rect 2700 5120 2964 5148
rect 2958 5108 2964 5120
rect 3016 5108 3022 5160
rect 3050 5108 3056 5160
rect 3108 5108 3114 5160
rect 5169 5151 5227 5157
rect 5169 5117 5181 5151
rect 5215 5148 5227 5151
rect 5258 5148 5264 5160
rect 5215 5120 5264 5148
rect 5215 5117 5227 5120
rect 5169 5111 5227 5117
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 5368 5080 5396 5188
rect 5445 5185 5457 5188
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 5552 5092 5580 5256
rect 6089 5253 6101 5256
rect 6135 5284 6147 5287
rect 6454 5284 6460 5296
rect 6135 5256 6460 5284
rect 6135 5253 6147 5256
rect 6089 5247 6147 5253
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 6914 5244 6920 5296
rect 6972 5244 6978 5296
rect 7466 5244 7472 5296
rect 7524 5284 7530 5296
rect 7524 5256 8064 5284
rect 7524 5244 7530 5256
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5185 5687 5219
rect 5629 5179 5687 5185
rect 5644 5148 5672 5179
rect 6546 5176 6552 5228
rect 6604 5216 6610 5228
rect 7662 5219 7720 5225
rect 7662 5216 7674 5219
rect 6604 5188 7674 5216
rect 6604 5176 6610 5188
rect 7662 5185 7674 5188
rect 7708 5185 7720 5219
rect 7662 5179 7720 5185
rect 5902 5148 5908 5160
rect 5644 5120 5908 5148
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 5442 5080 5448 5092
rect 2884 5052 4292 5080
rect 5368 5052 5448 5080
rect 2884 5024 2912 5052
rect 1578 4972 1584 5024
rect 1636 5012 1642 5024
rect 1765 5015 1823 5021
rect 1765 5012 1777 5015
rect 1636 4984 1777 5012
rect 1636 4972 1642 4984
rect 1765 4981 1777 4984
rect 1811 4981 1823 5015
rect 1765 4975 1823 4981
rect 2866 4972 2872 5024
rect 2924 4972 2930 5024
rect 3234 4972 3240 5024
rect 3292 5012 3298 5024
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3292 4984 3801 5012
rect 3292 4972 3298 4984
rect 3789 4981 3801 4984
rect 3835 5012 3847 5015
rect 4062 5012 4068 5024
rect 3835 4984 4068 5012
rect 3835 4981 3847 4984
rect 3789 4975 3847 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4264 5012 4292 5052
rect 5442 5040 5448 5052
rect 5500 5040 5506 5092
rect 5534 5040 5540 5092
rect 5592 5040 5598 5092
rect 6914 5080 6920 5092
rect 5644 5052 6920 5080
rect 5644 5012 5672 5052
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 4264 4984 5672 5012
rect 5905 5015 5963 5021
rect 5905 4981 5917 5015
rect 5951 5012 5963 5015
rect 6270 5012 6276 5024
rect 5951 4984 6276 5012
rect 5951 4981 5963 4984
rect 5905 4975 5963 4981
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 6549 5015 6607 5021
rect 6549 5012 6561 5015
rect 6512 4984 6561 5012
rect 6512 4972 6518 4984
rect 6549 4981 6561 4984
rect 6595 4981 6607 5015
rect 6549 4975 6607 4981
rect 7282 4972 7288 5024
rect 7340 5012 7346 5024
rect 7944 5012 7972 5111
rect 8036 5089 8064 5256
rect 8680 5256 9720 5284
rect 8202 5176 8208 5228
rect 8260 5176 8266 5228
rect 8680 5160 8708 5256
rect 9398 5176 9404 5228
rect 9456 5225 9462 5228
rect 9692 5225 9720 5256
rect 10318 5244 10324 5296
rect 10376 5244 10382 5296
rect 9456 5216 9468 5225
rect 9677 5219 9735 5225
rect 9456 5188 9501 5216
rect 9456 5179 9468 5188
rect 9677 5185 9689 5219
rect 9723 5185 9735 5219
rect 9677 5179 9735 5185
rect 9456 5176 9462 5179
rect 8662 5148 8668 5160
rect 8128 5120 8668 5148
rect 8021 5083 8079 5089
rect 8021 5049 8033 5083
rect 8067 5049 8079 5083
rect 8021 5043 8079 5049
rect 8128 5012 8156 5120
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 8220 5052 8432 5080
rect 8220 5024 8248 5052
rect 7340 4984 8156 5012
rect 7340 4972 7346 4984
rect 8202 4972 8208 5024
rect 8260 4972 8266 5024
rect 8294 4972 8300 5024
rect 8352 4972 8358 5024
rect 8404 5012 8432 5052
rect 9876 5052 10180 5080
rect 9876 5012 9904 5052
rect 8404 4984 9904 5012
rect 9950 4972 9956 5024
rect 10008 4972 10014 5024
rect 10152 5021 10180 5052
rect 10137 5015 10195 5021
rect 10137 4981 10149 5015
rect 10183 4981 10195 5015
rect 10137 4975 10195 4981
rect 1104 4922 10764 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 10764 4922
rect 1104 4848 10764 4870
rect 2866 4768 2872 4820
rect 2924 4768 2930 4820
rect 3053 4811 3111 4817
rect 3053 4777 3065 4811
rect 3099 4808 3111 4811
rect 4154 4808 4160 4820
rect 3099 4780 4160 4808
rect 3099 4777 3111 4780
rect 3053 4771 3111 4777
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 4341 4811 4399 4817
rect 4341 4808 4353 4811
rect 4304 4780 4353 4808
rect 4304 4768 4310 4780
rect 4341 4777 4353 4780
rect 4387 4777 4399 4811
rect 4341 4771 4399 4777
rect 5077 4811 5135 4817
rect 5077 4777 5089 4811
rect 5123 4777 5135 4811
rect 5077 4771 5135 4777
rect 3786 4700 3792 4752
rect 3844 4700 3850 4752
rect 5092 4740 5120 4771
rect 5166 4768 5172 4820
rect 5224 4808 5230 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 5224 4780 5273 4808
rect 5224 4768 5230 4780
rect 5261 4777 5273 4780
rect 5307 4777 5319 4811
rect 5261 4771 5319 4777
rect 6273 4811 6331 4817
rect 6273 4777 6285 4811
rect 6319 4808 6331 4811
rect 7374 4808 7380 4820
rect 6319 4780 7380 4808
rect 6319 4777 6331 4780
rect 6273 4771 6331 4777
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 8018 4768 8024 4820
rect 8076 4768 8082 4820
rect 8294 4768 8300 4820
rect 8352 4808 8358 4820
rect 10502 4808 10508 4820
rect 8352 4780 10508 4808
rect 8352 4768 8358 4780
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 5092 4712 6592 4740
rect 3510 4632 3516 4684
rect 3568 4632 3574 4684
rect 3804 4672 3832 4700
rect 3804 4644 6132 4672
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 3329 4607 3387 4613
rect 2639 4576 3188 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 3160 4480 3188 4576
rect 3329 4573 3341 4607
rect 3375 4604 3387 4607
rect 3970 4604 3976 4616
rect 3375 4576 3976 4604
rect 3375 4573 3387 4576
rect 3329 4567 3387 4573
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 4062 4564 4068 4616
rect 4120 4604 4126 4616
rect 4249 4607 4307 4613
rect 4249 4604 4261 4607
rect 4120 4576 4261 4604
rect 4120 4564 4126 4576
rect 4249 4573 4261 4576
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4479 4576 5304 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 3418 4496 3424 4548
rect 3476 4536 3482 4548
rect 4448 4536 4476 4567
rect 4890 4536 4896 4548
rect 3476 4508 4476 4536
rect 4832 4508 4896 4536
rect 3476 4496 3482 4508
rect 3142 4428 3148 4480
rect 3200 4428 3206 4480
rect 4430 4428 4436 4480
rect 4488 4468 4494 4480
rect 4832 4468 4860 4508
rect 4890 4496 4896 4508
rect 4948 4496 4954 4548
rect 5074 4496 5080 4548
rect 5132 4545 5138 4548
rect 5132 4539 5151 4545
rect 5139 4505 5151 4539
rect 5132 4499 5151 4505
rect 5132 4496 5138 4499
rect 4488 4440 4860 4468
rect 5276 4468 5304 4576
rect 5350 4564 5356 4616
rect 5408 4564 5414 4616
rect 6104 4613 6132 4644
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 5368 4536 5396 4564
rect 6380 4536 6408 4567
rect 5368 4508 6408 4536
rect 6454 4496 6460 4548
rect 6512 4496 6518 4548
rect 6564 4536 6592 4712
rect 9858 4632 9864 4684
rect 9916 4632 9922 4684
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4604 6699 4607
rect 7282 4604 7288 4616
rect 6687 4576 7288 4604
rect 6687 4573 6699 4576
rect 6641 4567 6699 4573
rect 7282 4564 7288 4576
rect 7340 4564 7346 4616
rect 9876 4604 9904 4632
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 7852 4576 10241 4604
rect 6914 4545 6920 4548
rect 6886 4539 6920 4545
rect 6564 4508 6776 4536
rect 6472 4468 6500 4496
rect 5276 4440 6500 4468
rect 4488 4428 4494 4440
rect 6546 4428 6552 4480
rect 6604 4428 6610 4480
rect 6748 4468 6776 4508
rect 6886 4505 6898 4539
rect 6886 4499 6920 4505
rect 6914 4496 6920 4499
rect 6972 4496 6978 4548
rect 7006 4496 7012 4548
rect 7064 4536 7070 4548
rect 7852 4536 7880 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 9858 4536 9864 4548
rect 7064 4508 7880 4536
rect 7944 4508 9864 4536
rect 7064 4496 7070 4508
rect 7944 4468 7972 4508
rect 9858 4496 9864 4508
rect 9916 4496 9922 4548
rect 6748 4440 7972 4468
rect 10410 4428 10416 4480
rect 10468 4428 10474 4480
rect 1104 4378 10764 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 10764 4378
rect 1104 4304 10764 4326
rect 1486 4224 1492 4276
rect 1544 4224 1550 4276
rect 2218 4267 2276 4273
rect 2218 4264 2230 4267
rect 1688 4236 2230 4264
rect 1504 4196 1532 4224
rect 1581 4199 1639 4205
rect 1581 4196 1593 4199
rect 1504 4168 1593 4196
rect 1581 4165 1593 4168
rect 1627 4165 1639 4199
rect 1581 4159 1639 4165
rect 1210 4088 1216 4140
rect 1268 4128 1274 4140
rect 1688 4128 1716 4236
rect 2218 4233 2230 4236
rect 2264 4233 2276 4267
rect 2218 4227 2276 4233
rect 2777 4267 2835 4273
rect 2777 4233 2789 4267
rect 2823 4264 2835 4267
rect 3142 4264 3148 4276
rect 2823 4236 3148 4264
rect 2823 4233 2835 4236
rect 2777 4227 2835 4233
rect 3142 4224 3148 4236
rect 3200 4264 3206 4276
rect 5994 4264 6000 4276
rect 3200 4236 6000 4264
rect 3200 4224 3206 4236
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 6546 4224 6552 4276
rect 6604 4264 6610 4276
rect 9674 4264 9680 4276
rect 6604 4236 9680 4264
rect 6604 4224 6610 4236
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 2406 4156 2412 4208
rect 2464 4156 2470 4208
rect 2593 4199 2651 4205
rect 2593 4165 2605 4199
rect 2639 4196 2651 4199
rect 3050 4196 3056 4208
rect 2639 4168 3056 4196
rect 2639 4165 2651 4168
rect 2593 4159 2651 4165
rect 3050 4156 3056 4168
rect 3108 4156 3114 4208
rect 6086 4156 6092 4208
rect 6144 4196 6150 4208
rect 6144 4168 6592 4196
rect 6144 4156 6150 4168
rect 1268 4100 1716 4128
rect 1765 4131 1823 4137
rect 1268 4088 1274 4100
rect 1765 4097 1777 4131
rect 1811 4097 1823 4131
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 1765 4091 1823 4097
rect 1872 4100 2053 4128
rect 1394 4020 1400 4072
rect 1452 4060 1458 4072
rect 1780 4060 1808 4091
rect 1872 4072 1900 4100
rect 2041 4097 2053 4100
rect 2087 4097 2099 4131
rect 2041 4091 2099 4097
rect 2130 4088 2136 4140
rect 2188 4088 2194 4140
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4128 2375 4131
rect 2498 4128 2504 4140
rect 2363 4100 2504 4128
rect 2363 4097 2375 4100
rect 2317 4091 2375 4097
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2958 4128 2964 4140
rect 2731 4100 2964 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 3344 4100 4936 4128
rect 3344 4072 3372 4100
rect 1452 4032 1808 4060
rect 1452 4020 1458 4032
rect 1854 4020 1860 4072
rect 1912 4060 1918 4072
rect 1912 4032 2084 4060
rect 1912 4020 1918 4032
rect 1762 3952 1768 4004
rect 1820 3992 1826 4004
rect 1949 3995 2007 4001
rect 1949 3992 1961 3995
rect 1820 3964 1961 3992
rect 1820 3952 1826 3964
rect 1949 3961 1961 3964
rect 1995 3961 2007 3995
rect 2056 3992 2084 4032
rect 2332 4032 2544 4060
rect 2332 3992 2360 4032
rect 2056 3964 2360 3992
rect 2516 3992 2544 4032
rect 2590 4020 2596 4072
rect 2648 4060 2654 4072
rect 3326 4060 3332 4072
rect 2648 4032 3332 4060
rect 2648 4020 2654 4032
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 4522 4020 4528 4072
rect 4580 4060 4586 4072
rect 4801 4063 4859 4069
rect 4801 4060 4813 4063
rect 4580 4032 4813 4060
rect 4580 4020 4586 4032
rect 4801 4029 4813 4032
rect 4847 4029 4859 4063
rect 4908 4060 4936 4100
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 5534 4128 5540 4140
rect 5040 4100 5540 4128
rect 5040 4088 5046 4100
rect 5534 4088 5540 4100
rect 5592 4128 5598 4140
rect 6178 4128 6184 4140
rect 5592 4100 6184 4128
rect 5592 4088 5598 4100
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 5074 4060 5080 4072
rect 4908 4032 5080 4060
rect 4801 4023 4859 4029
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 5169 4063 5227 4069
rect 5169 4029 5181 4063
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 5261 4063 5319 4069
rect 5261 4029 5273 4063
rect 5307 4060 5319 4063
rect 5350 4060 5356 4072
rect 5307 4032 5356 4060
rect 5307 4029 5319 4032
rect 5261 4023 5319 4029
rect 4614 3992 4620 4004
rect 2516 3964 4620 3992
rect 1949 3955 2007 3961
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 4706 3952 4712 4004
rect 4764 3992 4770 4004
rect 5184 3992 5212 4023
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 6454 4060 6460 4072
rect 5460 4032 6460 4060
rect 5460 3992 5488 4032
rect 6454 4020 6460 4032
rect 6512 4020 6518 4072
rect 6564 4060 6592 4168
rect 6638 4156 6644 4208
rect 6696 4156 6702 4208
rect 6822 4156 6828 4208
rect 6880 4156 6886 4208
rect 7025 4199 7083 4205
rect 7025 4196 7037 4199
rect 6932 4168 7037 4196
rect 6656 4128 6684 4156
rect 6932 4128 6960 4168
rect 7025 4165 7037 4168
rect 7071 4165 7083 4199
rect 7621 4199 7679 4205
rect 7621 4196 7633 4199
rect 7025 4159 7083 4165
rect 7116 4168 7633 4196
rect 6656 4100 6960 4128
rect 7116 4060 7144 4168
rect 7621 4165 7633 4168
rect 7667 4165 7679 4199
rect 7621 4159 7679 4165
rect 7834 4156 7840 4208
rect 7892 4156 7898 4208
rect 8570 4156 8576 4208
rect 8628 4156 8634 4208
rect 8588 4128 8616 4156
rect 6564 4032 7144 4060
rect 7208 4100 8616 4128
rect 5810 3992 5816 4004
rect 4764 3964 5488 3992
rect 5552 3964 5816 3992
rect 4764 3952 4770 3964
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 2130 3924 2136 3936
rect 1636 3896 2136 3924
rect 1636 3884 1642 3896
rect 2130 3884 2136 3896
rect 2188 3924 2194 3936
rect 2590 3924 2596 3936
rect 2188 3896 2596 3924
rect 2188 3884 2194 3896
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 2682 3884 2688 3936
rect 2740 3924 2746 3936
rect 2961 3927 3019 3933
rect 2961 3924 2973 3927
rect 2740 3896 2973 3924
rect 2740 3884 2746 3896
rect 2961 3893 2973 3896
rect 3007 3893 3019 3927
rect 2961 3887 3019 3893
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 5552 3924 5580 3964
rect 5810 3952 5816 3964
rect 5868 3992 5874 4004
rect 7208 4001 7236 4100
rect 7193 3995 7251 4001
rect 5868 3964 7144 3992
rect 5868 3952 5874 3964
rect 3844 3896 5580 3924
rect 3844 3884 3850 3896
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 7009 3927 7067 3933
rect 7009 3924 7021 3927
rect 5960 3896 7021 3924
rect 5960 3884 5966 3896
rect 7009 3893 7021 3896
rect 7055 3893 7067 3927
rect 7116 3924 7144 3964
rect 7193 3961 7205 3995
rect 7239 3961 7251 3995
rect 7193 3955 7251 3961
rect 7374 3952 7380 4004
rect 7432 3992 7438 4004
rect 7432 3964 9674 3992
rect 7432 3952 7438 3964
rect 7469 3927 7527 3933
rect 7469 3924 7481 3927
rect 7116 3896 7481 3924
rect 7009 3887 7067 3893
rect 7469 3893 7481 3896
rect 7515 3893 7527 3927
rect 7469 3887 7527 3893
rect 7653 3927 7711 3933
rect 7653 3893 7665 3927
rect 7699 3924 7711 3927
rect 8938 3924 8944 3936
rect 7699 3896 8944 3924
rect 7699 3893 7711 3896
rect 7653 3887 7711 3893
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9646 3924 9674 3964
rect 10042 3924 10048 3936
rect 9646 3896 10048 3924
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 1104 3834 10764 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 10764 3834
rect 1104 3760 10764 3782
rect 4798 3680 4804 3732
rect 4856 3680 4862 3732
rect 7009 3723 7067 3729
rect 5644 3692 6960 3720
rect 5644 3652 5672 3692
rect 2148 3624 5672 3652
rect 2038 3544 2044 3596
rect 2096 3544 2102 3596
rect 2148 3525 2176 3624
rect 3602 3544 3608 3596
rect 3660 3544 3666 3596
rect 5258 3584 5264 3596
rect 4908 3556 5264 3584
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3516 3019 3519
rect 3620 3516 3648 3544
rect 4908 3528 4936 3556
rect 5258 3544 5264 3556
rect 5316 3584 5322 3596
rect 5629 3587 5687 3593
rect 5629 3584 5641 3587
rect 5316 3556 5641 3584
rect 5316 3544 5322 3556
rect 5629 3553 5641 3556
rect 5675 3553 5687 3587
rect 6932 3584 6960 3692
rect 7009 3689 7021 3723
rect 7055 3720 7067 3723
rect 8478 3720 8484 3732
rect 7055 3692 8484 3720
rect 7055 3689 7067 3692
rect 7009 3683 7067 3689
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 9766 3720 9772 3732
rect 8772 3692 9772 3720
rect 7190 3612 7196 3664
rect 7248 3612 7254 3664
rect 7374 3612 7380 3664
rect 7432 3612 7438 3664
rect 8294 3652 8300 3664
rect 7576 3624 8300 3652
rect 7576 3584 7604 3624
rect 8294 3612 8300 3624
rect 8352 3612 8358 3664
rect 6932 3556 7604 3584
rect 7653 3587 7711 3593
rect 5629 3547 5687 3553
rect 7653 3553 7665 3587
rect 7699 3584 7711 3587
rect 8110 3584 8116 3596
rect 7699 3556 8116 3584
rect 7699 3553 7711 3556
rect 7653 3547 7711 3553
rect 8110 3544 8116 3556
rect 8168 3584 8174 3596
rect 8772 3584 8800 3692
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 9858 3680 9864 3732
rect 9916 3680 9922 3732
rect 9309 3655 9367 3661
rect 9309 3621 9321 3655
rect 9355 3652 9367 3655
rect 9355 3624 9812 3652
rect 9355 3621 9367 3624
rect 9309 3615 9367 3621
rect 8168 3556 8800 3584
rect 8168 3544 8174 3556
rect 9784 3528 9812 3624
rect 3007 3488 3648 3516
rect 4709 3519 4767 3525
rect 3007 3485 3019 3488
rect 2961 3479 3019 3485
rect 4709 3485 4721 3519
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 2406 3408 2412 3460
rect 2464 3448 2470 3460
rect 2682 3448 2688 3460
rect 2464 3420 2688 3448
rect 2464 3408 2470 3420
rect 2682 3408 2688 3420
rect 2740 3448 2746 3460
rect 4724 3448 4752 3479
rect 4890 3476 4896 3528
rect 4948 3476 4954 3528
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3485 5043 3519
rect 4985 3479 5043 3485
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5442 3516 5448 3528
rect 5215 3488 5448 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 2740 3420 4752 3448
rect 5000 3448 5028 3479
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 5534 3476 5540 3528
rect 5592 3476 5598 3528
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 5885 3519 5943 3525
rect 5885 3516 5897 3519
rect 5776 3488 5897 3516
rect 5776 3476 5782 3488
rect 5885 3485 5897 3488
rect 5931 3485 5943 3519
rect 5885 3479 5943 3485
rect 6178 3476 6184 3528
rect 6236 3516 6242 3528
rect 9033 3519 9091 3525
rect 9033 3516 9045 3519
rect 6236 3488 9045 3516
rect 6236 3476 6242 3488
rect 9033 3485 9045 3488
rect 9079 3485 9091 3519
rect 9033 3479 9091 3485
rect 9490 3476 9496 3528
rect 9548 3476 9554 3528
rect 9766 3476 9772 3528
rect 9824 3476 9830 3528
rect 10134 3476 10140 3528
rect 10192 3476 10198 3528
rect 10226 3476 10232 3528
rect 10284 3516 10290 3528
rect 10778 3516 10784 3528
rect 10284 3488 10784 3516
rect 10284 3476 10290 3488
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 6362 3448 6368 3460
rect 5000 3420 6368 3448
rect 2740 3408 2746 3420
rect 6362 3408 6368 3420
rect 6420 3408 6426 3460
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 9309 3451 9367 3457
rect 9309 3448 9321 3451
rect 6512 3420 9321 3448
rect 6512 3408 6518 3420
rect 9309 3417 9321 3420
rect 9355 3417 9367 3451
rect 9309 3411 9367 3417
rect 9677 3451 9735 3457
rect 9677 3417 9689 3451
rect 9723 3448 9735 3451
rect 10152 3448 10180 3476
rect 10686 3448 10692 3460
rect 9723 3420 10180 3448
rect 10336 3420 10692 3448
rect 9723 3417 9735 3420
rect 9677 3411 9735 3417
rect 3145 3383 3203 3389
rect 3145 3349 3157 3383
rect 3191 3380 3203 3383
rect 6270 3380 6276 3392
rect 3191 3352 6276 3380
rect 3191 3349 3203 3352
rect 3145 3343 3203 3349
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 6638 3340 6644 3392
rect 6696 3380 6702 3392
rect 9125 3383 9183 3389
rect 9125 3380 9137 3383
rect 6696 3352 9137 3380
rect 6696 3340 6702 3352
rect 9125 3349 9137 3352
rect 9171 3380 9183 3383
rect 9214 3380 9220 3392
rect 9171 3352 9220 3380
rect 9171 3349 9183 3352
rect 9125 3343 9183 3349
rect 9214 3340 9220 3352
rect 9272 3340 9278 3392
rect 9324 3380 9352 3411
rect 10042 3380 10048 3392
rect 9324 3352 10048 3380
rect 10042 3340 10048 3352
rect 10100 3380 10106 3392
rect 10336 3380 10364 3420
rect 10686 3408 10692 3420
rect 10744 3408 10750 3460
rect 10100 3352 10364 3380
rect 10100 3340 10106 3352
rect 10410 3340 10416 3392
rect 10468 3340 10474 3392
rect 1104 3290 10764 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 10764 3290
rect 1104 3216 10764 3238
rect 2777 3179 2835 3185
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 4154 3176 4160 3188
rect 2823 3148 4160 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 4249 3179 4307 3185
rect 4249 3145 4261 3179
rect 4295 3176 4307 3179
rect 4982 3176 4988 3188
rect 4295 3148 4988 3176
rect 4295 3145 4307 3148
rect 4249 3139 4307 3145
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 5721 3179 5779 3185
rect 5721 3145 5733 3179
rect 5767 3176 5779 3179
rect 5810 3176 5816 3188
rect 5767 3148 5816 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 6549 3179 6607 3185
rect 6549 3145 6561 3179
rect 6595 3176 6607 3179
rect 6730 3176 6736 3188
rect 6595 3148 6736 3176
rect 6595 3145 6607 3148
rect 6549 3139 6607 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 7282 3176 7288 3188
rect 7024 3148 7288 3176
rect 4608 3111 4666 3117
rect 1412 3080 4476 3108
rect 1412 3049 1440 3080
rect 1670 3049 1676 3052
rect 1397 3043 1455 3049
rect 1397 3009 1409 3043
rect 1443 3009 1455 3043
rect 1664 3040 1676 3049
rect 1631 3012 1676 3040
rect 1397 3003 1455 3009
rect 1664 3003 1676 3012
rect 1670 3000 1676 3003
rect 1728 3000 1734 3052
rect 2958 3040 2964 3052
rect 2746 3012 2964 3040
rect 2498 2932 2504 2984
rect 2556 2972 2562 2984
rect 2746 2972 2774 3012
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3040 3111 3043
rect 3142 3040 3148 3052
rect 3099 3012 3148 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3040 3295 3043
rect 3786 3040 3792 3052
rect 3283 3012 3792 3040
rect 3283 3009 3295 3012
rect 3237 3003 3295 3009
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 3970 3040 3976 3052
rect 3927 3012 3976 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3040 4123 3043
rect 4448 3040 4476 3080
rect 4608 3077 4620 3111
rect 4654 3108 4666 3111
rect 4706 3108 4712 3120
rect 4654 3080 4712 3108
rect 4654 3077 4666 3080
rect 4608 3071 4666 3077
rect 4706 3068 4712 3080
rect 4764 3068 4770 3120
rect 5074 3068 5080 3120
rect 5132 3068 5138 3120
rect 5644 3080 6408 3108
rect 4890 3040 4896 3052
rect 4111 3012 4292 3040
rect 4111 3009 4123 3012
rect 4065 3003 4123 3009
rect 2556 2944 2774 2972
rect 2556 2932 2562 2944
rect 2869 2839 2927 2845
rect 2869 2805 2881 2839
rect 2915 2836 2927 2839
rect 4154 2836 4160 2848
rect 2915 2808 4160 2836
rect 2915 2805 2927 2808
rect 2869 2799 2927 2805
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 4264 2836 4292 3012
rect 4448 3012 4896 3040
rect 4341 2975 4399 2981
rect 4341 2941 4353 2975
rect 4387 2972 4399 2975
rect 4448 2972 4476 3012
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 5092 3040 5120 3068
rect 5644 3052 5672 3080
rect 5092 3012 5580 3040
rect 4387 2944 4476 2972
rect 5552 2972 5580 3012
rect 5626 3000 5632 3052
rect 5684 3000 5690 3052
rect 6270 3000 6276 3052
rect 6328 3000 6334 3052
rect 6380 3049 6408 3080
rect 7024 3049 7052 3148
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 9030 3176 9036 3188
rect 8435 3148 9036 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 9214 3136 9220 3188
rect 9272 3136 9278 3188
rect 9398 3136 9404 3188
rect 9456 3136 9462 3188
rect 9232 3108 9260 3136
rect 9232 3080 10180 3108
rect 10152 3052 10180 3080
rect 10870 3068 10876 3120
rect 10928 3068 10934 3120
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3009 7067 3043
rect 7265 3043 7323 3049
rect 7265 3040 7277 3043
rect 7009 3003 7067 3009
rect 7116 3012 7277 3040
rect 6288 2972 6316 3000
rect 7116 2972 7144 3012
rect 7265 3009 7277 3012
rect 7311 3009 7323 3043
rect 7265 3003 7323 3009
rect 9122 3000 9128 3052
rect 9180 3040 9186 3052
rect 9401 3043 9459 3049
rect 9401 3040 9413 3043
rect 9180 3012 9413 3040
rect 9180 3000 9186 3012
rect 9401 3009 9413 3012
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 9766 3000 9772 3052
rect 9824 3000 9830 3052
rect 10042 3000 10048 3052
rect 10100 3000 10106 3052
rect 10134 3000 10140 3052
rect 10192 3000 10198 3052
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10888 3040 10916 3068
rect 10376 3012 10916 3040
rect 10376 3000 10382 3012
rect 5552 2944 6224 2972
rect 6288 2944 7144 2972
rect 4387 2941 4399 2944
rect 4341 2935 4399 2941
rect 5350 2864 5356 2916
rect 5408 2904 5414 2916
rect 6196 2904 6224 2944
rect 10226 2932 10232 2984
rect 10284 2932 10290 2984
rect 6638 2904 6644 2916
rect 5408 2876 5856 2904
rect 6196 2876 6644 2904
rect 5408 2864 5414 2876
rect 5718 2836 5724 2848
rect 4264 2808 5724 2836
rect 5718 2796 5724 2808
rect 5776 2796 5782 2848
rect 5828 2836 5856 2876
rect 6638 2864 6644 2876
rect 6696 2864 6702 2916
rect 10244 2836 10272 2932
rect 5828 2808 10272 2836
rect 1104 2746 10764 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 10764 2746
rect 1104 2672 10764 2694
rect 934 2592 940 2644
rect 992 2632 998 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 992 2604 2421 2632
rect 992 2592 998 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 5353 2635 5411 2641
rect 2409 2595 2467 2601
rect 2516 2604 2774 2632
rect 2516 2573 2544 2604
rect 2501 2567 2559 2573
rect 2501 2533 2513 2567
rect 2547 2533 2559 2567
rect 2501 2527 2559 2533
rect 750 2456 756 2508
rect 808 2456 814 2508
rect 1854 2456 1860 2508
rect 1912 2496 1918 2508
rect 2133 2499 2191 2505
rect 2133 2496 2145 2499
rect 1912 2468 2145 2496
rect 1912 2456 1918 2468
rect 2133 2465 2145 2468
rect 2179 2465 2191 2499
rect 2133 2459 2191 2465
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2496 2283 2499
rect 2590 2496 2596 2508
rect 2271 2468 2596 2496
rect 2271 2465 2283 2468
rect 2225 2459 2283 2465
rect 2590 2456 2596 2468
rect 2648 2456 2654 2508
rect 2746 2496 2774 2604
rect 5353 2601 5365 2635
rect 5399 2632 5411 2635
rect 6730 2632 6736 2644
rect 5399 2604 6736 2632
rect 5399 2601 5411 2604
rect 5353 2595 5411 2601
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 6822 2592 6828 2644
rect 6880 2592 6886 2644
rect 4430 2524 4436 2576
rect 4488 2564 4494 2576
rect 4985 2567 5043 2573
rect 4985 2564 4997 2567
rect 4488 2536 4997 2564
rect 4488 2524 4494 2536
rect 4985 2533 4997 2536
rect 5031 2533 5043 2567
rect 4985 2527 5043 2533
rect 5626 2524 5632 2576
rect 5684 2564 5690 2576
rect 6089 2567 6147 2573
rect 6089 2564 6101 2567
rect 5684 2536 6101 2564
rect 5684 2524 5690 2536
rect 6089 2533 6101 2536
rect 6135 2533 6147 2567
rect 6089 2527 6147 2533
rect 6840 2496 6868 2592
rect 2746 2468 6868 2496
rect 768 2428 796 2456
rect 1949 2431 2007 2437
rect 1949 2428 1961 2431
rect 768 2400 1961 2428
rect 1688 2292 1716 2400
rect 1949 2397 1961 2400
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 1762 2320 1768 2372
rect 1820 2360 1826 2372
rect 2056 2360 2084 2391
rect 2314 2388 2320 2440
rect 2372 2428 2378 2440
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2372 2400 2513 2428
rect 2372 2388 2378 2400
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2428 6147 2431
rect 7374 2428 7380 2440
rect 6135 2400 7380 2428
rect 6135 2397 6147 2400
rect 6089 2391 6147 2397
rect 1820 2332 2084 2360
rect 1820 2320 1826 2332
rect 2406 2320 2412 2372
rect 2464 2360 2470 2372
rect 2700 2360 2728 2391
rect 2464 2332 2728 2360
rect 2464 2320 2470 2332
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 5353 2363 5411 2369
rect 5353 2360 5365 2363
rect 4212 2332 5365 2360
rect 4212 2320 4218 2332
rect 5353 2329 5365 2332
rect 5399 2329 5411 2363
rect 5920 2360 5948 2391
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 8110 2388 8116 2440
rect 8168 2388 8174 2440
rect 8202 2388 8208 2440
rect 8260 2388 8266 2440
rect 9950 2388 9956 2440
rect 10008 2388 10014 2440
rect 10226 2388 10232 2440
rect 10284 2388 10290 2440
rect 8128 2360 8156 2388
rect 5353 2323 5411 2329
rect 5460 2332 8156 2360
rect 5460 2292 5488 2332
rect 1688 2264 5488 2292
rect 5537 2295 5595 2301
rect 5537 2261 5549 2295
rect 5583 2292 5595 2295
rect 8220 2292 8248 2388
rect 5583 2264 8248 2292
rect 5583 2261 5595 2264
rect 5537 2255 5595 2261
rect 10134 2252 10140 2304
rect 10192 2252 10198 2304
rect 10413 2295 10471 2301
rect 10413 2261 10425 2295
rect 10459 2292 10471 2295
rect 10459 2264 10916 2292
rect 10459 2261 10471 2264
rect 10413 2255 10471 2261
rect 10888 2236 10916 2264
rect 1104 2202 10764 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 10764 2202
rect 10870 2184 10876 2236
rect 10928 2184 10934 2236
rect 1104 2128 10764 2150
rect 750 2048 756 2100
rect 808 2088 814 2100
rect 7282 2088 7288 2100
rect 808 2060 7288 2088
rect 808 2048 814 2060
rect 7282 2048 7288 2060
rect 7340 2048 7346 2100
<< via1 >>
rect 1676 11568 1728 11620
rect 8576 11568 8628 11620
rect 2596 11500 2648 11552
rect 4528 11500 4580 11552
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 6950 11398 7002 11450
rect 7014 11398 7066 11450
rect 7078 11398 7130 11450
rect 7142 11398 7194 11450
rect 7206 11398 7258 11450
rect 1676 11296 1728 11348
rect 3424 11296 3476 11348
rect 1768 11228 1820 11280
rect 1584 11160 1636 11212
rect 2596 11203 2648 11212
rect 2596 11169 2605 11203
rect 2605 11169 2639 11203
rect 2639 11169 2648 11203
rect 2596 11160 2648 11169
rect 3056 11228 3108 11280
rect 3148 11228 3200 11280
rect 3700 11228 3752 11280
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 1860 11092 1912 11144
rect 2504 11024 2556 11076
rect 4160 11160 4212 11212
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 5632 11228 5684 11280
rect 8392 11228 8444 11280
rect 9680 11296 9732 11348
rect 8760 11271 8812 11280
rect 8760 11237 8769 11271
rect 8769 11237 8803 11271
rect 8803 11237 8812 11271
rect 8760 11228 8812 11237
rect 3056 11067 3108 11076
rect 3056 11033 3065 11067
rect 3065 11033 3099 11067
rect 3099 11033 3108 11067
rect 3056 11024 3108 11033
rect 3700 11024 3752 11076
rect 3792 11024 3844 11076
rect 5724 11135 5776 11144
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 5816 11135 5868 11144
rect 5816 11101 5825 11135
rect 5825 11101 5859 11135
rect 5859 11101 5868 11135
rect 5816 11092 5868 11101
rect 8484 11092 8536 11144
rect 4620 11067 4672 11076
rect 4620 11033 4629 11067
rect 4629 11033 4663 11067
rect 4663 11033 4672 11067
rect 4620 11024 4672 11033
rect 5540 11067 5592 11076
rect 5540 11033 5549 11067
rect 5549 11033 5583 11067
rect 5583 11033 5592 11067
rect 5540 11024 5592 11033
rect 7472 11024 7524 11076
rect 9404 11024 9456 11076
rect 3516 10999 3568 11008
rect 3516 10965 3525 10999
rect 3525 10965 3559 10999
rect 3559 10965 3568 10999
rect 3516 10956 3568 10965
rect 4528 10956 4580 11008
rect 5724 10956 5776 11008
rect 7196 10956 7248 11008
rect 10048 10956 10100 11008
rect 2610 10854 2662 10906
rect 2674 10854 2726 10906
rect 2738 10854 2790 10906
rect 2802 10854 2854 10906
rect 2866 10854 2918 10906
rect 7610 10854 7662 10906
rect 7674 10854 7726 10906
rect 7738 10854 7790 10906
rect 7802 10854 7854 10906
rect 7866 10854 7918 10906
rect 1768 10752 1820 10804
rect 1860 10795 1912 10804
rect 1860 10761 1869 10795
rect 1869 10761 1903 10795
rect 1903 10761 1912 10795
rect 1860 10752 1912 10761
rect 3148 10752 3200 10804
rect 4068 10752 4120 10804
rect 7196 10795 7248 10804
rect 7196 10761 7205 10795
rect 7205 10761 7239 10795
rect 7239 10761 7248 10795
rect 7196 10752 7248 10761
rect 7932 10752 7984 10804
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 1676 10616 1728 10668
rect 4160 10684 4212 10736
rect 4620 10684 4672 10736
rect 5632 10684 5684 10736
rect 9588 10752 9640 10804
rect 2504 10548 2556 10600
rect 3056 10659 3108 10668
rect 3056 10625 3065 10659
rect 3065 10625 3099 10659
rect 3099 10625 3108 10659
rect 3056 10616 3108 10625
rect 3240 10616 3292 10668
rect 3884 10616 3936 10668
rect 5816 10616 5868 10668
rect 7656 10616 7708 10668
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 9404 10684 9456 10736
rect 3792 10548 3844 10600
rect 1860 10412 1912 10464
rect 2320 10455 2372 10464
rect 2320 10421 2329 10455
rect 2329 10421 2363 10455
rect 2363 10421 2372 10455
rect 2320 10412 2372 10421
rect 6000 10480 6052 10532
rect 6368 10480 6420 10532
rect 8024 10548 8076 10600
rect 8300 10659 8352 10668
rect 8300 10625 8309 10659
rect 8309 10625 8343 10659
rect 8343 10625 8352 10659
rect 8300 10616 8352 10625
rect 8392 10616 8444 10668
rect 8668 10616 8720 10668
rect 8208 10480 8260 10532
rect 8484 10480 8536 10532
rect 3516 10412 3568 10464
rect 3700 10412 3752 10464
rect 6460 10412 6512 10464
rect 8852 10412 8904 10464
rect 8944 10455 8996 10464
rect 8944 10421 8953 10455
rect 8953 10421 8987 10455
rect 8987 10421 8996 10455
rect 8944 10412 8996 10421
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 6950 10310 7002 10362
rect 7014 10310 7066 10362
rect 7078 10310 7130 10362
rect 7142 10310 7194 10362
rect 7206 10310 7258 10362
rect 2872 10208 2924 10260
rect 3976 10208 4028 10260
rect 4528 10251 4580 10260
rect 4528 10217 4537 10251
rect 4537 10217 4571 10251
rect 4571 10217 4580 10251
rect 4528 10208 4580 10217
rect 7840 10208 7892 10260
rect 7932 10208 7984 10260
rect 8484 10208 8536 10260
rect 8576 10208 8628 10260
rect 9864 10208 9916 10260
rect 10876 10208 10928 10260
rect 6276 10140 6328 10192
rect 3608 10115 3660 10124
rect 3608 10081 3617 10115
rect 3617 10081 3651 10115
rect 3651 10081 3660 10115
rect 3608 10072 3660 10081
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2964 10004 3016 10056
rect 3148 10004 3200 10056
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 3700 10004 3752 10056
rect 940 9936 992 9988
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 4620 10004 4672 10056
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 6092 10072 6144 10124
rect 6184 10004 6236 10056
rect 7656 10072 7708 10124
rect 8300 10072 8352 10124
rect 6644 10004 6696 10056
rect 8024 10004 8076 10056
rect 9036 10004 9088 10056
rect 9128 10004 9180 10056
rect 4712 9936 4764 9988
rect 6920 9936 6972 9988
rect 1676 9868 1728 9920
rect 2504 9868 2556 9920
rect 2872 9868 2924 9920
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 3332 9868 3384 9920
rect 4252 9911 4304 9920
rect 4252 9877 4261 9911
rect 4261 9877 4295 9911
rect 4295 9877 4304 9911
rect 4252 9868 4304 9877
rect 4436 9868 4488 9920
rect 4896 9911 4948 9920
rect 4896 9877 4905 9911
rect 4905 9877 4939 9911
rect 4939 9877 4948 9911
rect 4896 9868 4948 9877
rect 6092 9911 6144 9920
rect 6092 9877 6101 9911
rect 6101 9877 6135 9911
rect 6135 9877 6144 9911
rect 6092 9868 6144 9877
rect 7380 9868 7432 9920
rect 9772 9936 9824 9988
rect 9864 9979 9916 9988
rect 9864 9945 9873 9979
rect 9873 9945 9907 9979
rect 9907 9945 9916 9979
rect 9864 9936 9916 9945
rect 8300 9868 8352 9920
rect 9220 9868 9272 9920
rect 9588 9868 9640 9920
rect 10692 9868 10744 9920
rect 10784 9868 10836 9920
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 7610 9766 7662 9818
rect 7674 9766 7726 9818
rect 7738 9766 7790 9818
rect 7802 9766 7854 9818
rect 7866 9766 7918 9818
rect 4712 9664 4764 9716
rect 6000 9707 6052 9716
rect 6000 9673 6009 9707
rect 6009 9673 6043 9707
rect 6043 9673 6052 9707
rect 6000 9664 6052 9673
rect 7564 9664 7616 9716
rect 8024 9664 8076 9716
rect 4620 9596 4672 9648
rect 4896 9639 4948 9648
rect 4896 9605 4914 9639
rect 4914 9605 4948 9639
rect 4896 9596 4948 9605
rect 6644 9596 6696 9648
rect 664 9528 716 9580
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 4436 9528 4488 9580
rect 5080 9528 5132 9580
rect 3700 9460 3752 9512
rect 4068 9460 4120 9512
rect 2780 9324 2832 9376
rect 2964 9324 3016 9376
rect 4160 9392 4212 9444
rect 3976 9324 4028 9376
rect 4068 9324 4120 9376
rect 6000 9392 6052 9444
rect 6920 9528 6972 9580
rect 7656 9528 7708 9580
rect 8300 9596 8352 9648
rect 9220 9664 9272 9716
rect 10508 9664 10560 9716
rect 9128 9596 9180 9648
rect 8116 9528 8168 9580
rect 10324 9596 10376 9648
rect 9404 9460 9456 9512
rect 7840 9392 7892 9444
rect 5816 9324 5868 9376
rect 6828 9324 6880 9376
rect 8024 9367 8076 9376
rect 8024 9333 8033 9367
rect 8033 9333 8067 9367
rect 8067 9333 8076 9367
rect 8024 9324 8076 9333
rect 8208 9367 8260 9376
rect 8208 9333 8217 9367
rect 8217 9333 8251 9367
rect 8251 9333 8260 9367
rect 8208 9324 8260 9333
rect 8576 9435 8628 9444
rect 8576 9401 8585 9435
rect 8585 9401 8619 9435
rect 8619 9401 8628 9435
rect 8576 9392 8628 9401
rect 9220 9392 9272 9444
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 10048 9528 10100 9580
rect 9128 9324 9180 9376
rect 9680 9324 9732 9376
rect 9772 9324 9824 9376
rect 9864 9324 9916 9376
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 10416 9367 10468 9376
rect 10416 9333 10425 9367
rect 10425 9333 10459 9367
rect 10459 9333 10468 9367
rect 10416 9324 10468 9333
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 1216 9052 1268 9104
rect 4804 9052 4856 9104
rect 7656 9120 7708 9172
rect 8300 9120 8352 9172
rect 8392 9120 8444 9172
rect 9220 9163 9272 9172
rect 9220 9129 9229 9163
rect 9229 9129 9263 9163
rect 9263 9129 9272 9163
rect 9220 9120 9272 9129
rect 10048 9163 10100 9172
rect 10048 9129 10057 9163
rect 10057 9129 10091 9163
rect 10091 9129 10100 9163
rect 10048 9120 10100 9129
rect 2872 8984 2924 9036
rect 2320 8848 2372 8900
rect 3240 8984 3292 9036
rect 3424 8984 3476 9036
rect 5816 8984 5868 9036
rect 7288 8984 7340 9036
rect 5908 8916 5960 8968
rect 6644 8916 6696 8968
rect 6736 8916 6788 8968
rect 3424 8848 3476 8900
rect 4896 8848 4948 8900
rect 5080 8848 5132 8900
rect 4344 8780 4396 8832
rect 5356 8780 5408 8832
rect 5540 8848 5592 8900
rect 6920 8780 6972 8832
rect 8024 8959 8076 8968
rect 8024 8925 8033 8959
rect 8033 8925 8067 8959
rect 8067 8925 8076 8959
rect 8024 8916 8076 8925
rect 8300 8916 8352 8968
rect 9220 8916 9272 8968
rect 9588 8959 9640 8968
rect 9588 8925 9597 8959
rect 9597 8925 9631 8959
rect 9631 8925 9640 8959
rect 9588 8916 9640 8925
rect 9956 8916 10008 8968
rect 8116 8848 8168 8900
rect 10232 8891 10284 8900
rect 10232 8857 10241 8891
rect 10241 8857 10275 8891
rect 10275 8857 10284 8891
rect 10232 8848 10284 8857
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 9496 8823 9548 8832
rect 9496 8789 9505 8823
rect 9505 8789 9539 8823
rect 9539 8789 9548 8823
rect 9496 8780 9548 8789
rect 9864 8823 9916 8832
rect 9864 8789 9873 8823
rect 9873 8789 9907 8823
rect 9907 8789 9916 8823
rect 9864 8780 9916 8789
rect 10140 8780 10192 8832
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 7610 8678 7662 8730
rect 7674 8678 7726 8730
rect 7738 8678 7790 8730
rect 7802 8678 7854 8730
rect 7866 8678 7918 8730
rect 3424 8576 3476 8628
rect 3976 8576 4028 8628
rect 4252 8576 4304 8628
rect 5908 8576 5960 8628
rect 8484 8576 8536 8628
rect 8944 8576 8996 8628
rect 1124 8372 1176 8424
rect 4712 8508 4764 8560
rect 5172 8440 5224 8492
rect 6000 8440 6052 8492
rect 9128 8440 9180 8492
rect 9680 8440 9732 8492
rect 3148 8372 3200 8424
rect 4068 8372 4120 8424
rect 4344 8372 4396 8424
rect 4160 8304 4212 8356
rect 4528 8304 4580 8356
rect 4804 8279 4856 8288
rect 4804 8245 4813 8279
rect 4813 8245 4847 8279
rect 4847 8245 4856 8279
rect 4804 8236 4856 8245
rect 5448 8236 5500 8288
rect 5540 8279 5592 8288
rect 5540 8245 5549 8279
rect 5549 8245 5583 8279
rect 5583 8245 5592 8279
rect 5540 8236 5592 8245
rect 6920 8304 6972 8356
rect 8300 8304 8352 8356
rect 9404 8236 9456 8288
rect 9864 8347 9916 8356
rect 9864 8313 9873 8347
rect 9873 8313 9907 8347
rect 9907 8313 9916 8347
rect 9864 8304 9916 8313
rect 10048 8279 10100 8288
rect 10048 8245 10057 8279
rect 10057 8245 10091 8279
rect 10091 8245 10100 8279
rect 10048 8236 10100 8245
rect 10416 8236 10468 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 4896 8032 4948 8084
rect 5264 8032 5316 8084
rect 8760 8032 8812 8084
rect 1308 7896 1360 7948
rect 7288 7896 7340 7948
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 5356 7828 5408 7880
rect 6184 7828 6236 7880
rect 6552 7828 6604 7880
rect 6736 7828 6788 7880
rect 8300 7896 8352 7948
rect 8760 7896 8812 7948
rect 8944 8032 8996 8084
rect 8944 7896 8996 7948
rect 8668 7828 8720 7880
rect 4896 7760 4948 7812
rect 10416 7828 10468 7880
rect 6092 7760 6144 7812
rect 6644 7760 6696 7812
rect 6920 7760 6972 7812
rect 8300 7760 8352 7812
rect 10600 7760 10652 7812
rect 2964 7692 3016 7744
rect 3424 7692 3476 7744
rect 3700 7692 3752 7744
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 5632 7692 5684 7744
rect 8760 7692 8812 7744
rect 9220 7735 9272 7744
rect 9220 7701 9229 7735
rect 9229 7701 9263 7735
rect 9263 7701 9272 7735
rect 9220 7692 9272 7701
rect 10416 7735 10468 7744
rect 10416 7701 10425 7735
rect 10425 7701 10459 7735
rect 10459 7701 10468 7735
rect 10416 7692 10468 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 2504 7488 2556 7540
rect 3700 7488 3752 7540
rect 3976 7488 4028 7540
rect 5448 7488 5500 7540
rect 3056 7420 3108 7472
rect 5540 7420 5592 7472
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 2688 7352 2740 7404
rect 4160 7352 4212 7404
rect 7472 7488 7524 7540
rect 8208 7488 8260 7540
rect 8944 7488 8996 7540
rect 10324 7488 10376 7540
rect 7380 7420 7432 7472
rect 4068 7327 4120 7336
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 4068 7284 4120 7293
rect 6828 7352 6880 7404
rect 8300 7352 8352 7404
rect 10600 7352 10652 7404
rect 6000 7284 6052 7336
rect 9496 7284 9548 7336
rect 6644 7216 6696 7268
rect 8944 7216 8996 7268
rect 9312 7216 9364 7268
rect 756 7148 808 7200
rect 4620 7148 4672 7200
rect 5908 7148 5960 7200
rect 7564 7148 7616 7200
rect 8760 7148 8812 7200
rect 9404 7148 9456 7200
rect 10324 7259 10376 7268
rect 10324 7225 10333 7259
rect 10333 7225 10367 7259
rect 10367 7225 10376 7259
rect 10324 7216 10376 7225
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 2688 6944 2740 6996
rect 3792 6987 3844 6996
rect 3792 6953 3801 6987
rect 3801 6953 3835 6987
rect 3835 6953 3844 6987
rect 3792 6944 3844 6953
rect 2228 6876 2280 6928
rect 5540 6944 5592 6996
rect 6828 6944 6880 6996
rect 7380 6944 7432 6996
rect 8668 6944 8720 6996
rect 10048 6944 10100 6996
rect 2504 6808 2556 6860
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 1952 6604 2004 6656
rect 2688 6740 2740 6792
rect 3240 6808 3292 6860
rect 3884 6808 3936 6860
rect 2136 6604 2188 6656
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 2596 6604 2648 6656
rect 2780 6647 2832 6656
rect 2780 6613 2789 6647
rect 2789 6613 2823 6647
rect 2823 6613 2832 6647
rect 2780 6604 2832 6613
rect 3332 6740 3384 6792
rect 5908 6808 5960 6860
rect 6368 6808 6420 6860
rect 6644 6808 6696 6860
rect 7380 6808 7432 6860
rect 3240 6715 3292 6724
rect 3240 6681 3249 6715
rect 3249 6681 3283 6715
rect 3283 6681 3292 6715
rect 3240 6672 3292 6681
rect 5264 6740 5316 6792
rect 5724 6740 5776 6792
rect 6092 6740 6144 6792
rect 8208 6740 8260 6792
rect 8300 6740 8352 6792
rect 3424 6647 3476 6656
rect 3424 6613 3449 6647
rect 3449 6613 3476 6647
rect 3424 6604 3476 6613
rect 3700 6604 3752 6656
rect 5448 6672 5500 6724
rect 6552 6672 6604 6724
rect 9312 6740 9364 6792
rect 8944 6672 8996 6724
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 10140 6672 10192 6724
rect 9588 6647 9640 6656
rect 9588 6613 9597 6647
rect 9597 6613 9631 6647
rect 9631 6613 9640 6647
rect 9588 6604 9640 6613
rect 10416 6647 10468 6656
rect 10416 6613 10425 6647
rect 10425 6613 10459 6647
rect 10459 6613 10468 6647
rect 10416 6604 10468 6613
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 1492 6400 1544 6452
rect 1860 6400 1912 6452
rect 2228 6400 2280 6452
rect 1308 6264 1360 6316
rect 2688 6375 2740 6384
rect 2688 6341 2697 6375
rect 2697 6341 2731 6375
rect 2731 6341 2740 6375
rect 2688 6332 2740 6341
rect 2872 6375 2924 6384
rect 2872 6341 2913 6375
rect 2913 6341 2924 6375
rect 2872 6332 2924 6341
rect 4344 6332 4396 6384
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 5632 6400 5684 6452
rect 5540 6332 5592 6384
rect 6092 6332 6144 6384
rect 6460 6443 6512 6452
rect 6460 6409 6469 6443
rect 6469 6409 6503 6443
rect 6503 6409 6512 6443
rect 6460 6400 6512 6409
rect 6644 6400 6696 6452
rect 7932 6400 7984 6452
rect 8208 6400 8260 6452
rect 8668 6400 8720 6452
rect 8944 6443 8996 6452
rect 8944 6409 8953 6443
rect 8953 6409 8987 6443
rect 8987 6409 8996 6443
rect 8944 6400 8996 6409
rect 9128 6400 9180 6452
rect 6736 6332 6788 6384
rect 6920 6332 6972 6384
rect 7656 6332 7708 6384
rect 7748 6332 7800 6384
rect 3792 6196 3844 6248
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 4252 6196 4304 6248
rect 6460 6196 6512 6248
rect 7104 6239 7156 6248
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 8484 6196 8536 6248
rect 9036 6332 9088 6384
rect 9220 6332 9272 6384
rect 9772 6332 9824 6384
rect 10324 6400 10376 6452
rect 10232 6332 10284 6384
rect 9404 6196 9456 6248
rect 1492 6128 1544 6180
rect 2228 6060 2280 6112
rect 2412 6060 2464 6112
rect 3792 6060 3844 6112
rect 3884 6103 3936 6112
rect 3884 6069 3893 6103
rect 3893 6069 3927 6103
rect 3927 6069 3936 6103
rect 3884 6060 3936 6069
rect 4988 6060 5040 6112
rect 5632 6060 5684 6112
rect 5724 6060 5776 6112
rect 8576 6128 8628 6180
rect 8944 6060 8996 6112
rect 9404 6103 9456 6112
rect 9404 6069 9413 6103
rect 9413 6069 9447 6103
rect 9447 6069 9456 6103
rect 9404 6060 9456 6069
rect 9496 6060 9548 6112
rect 10324 6060 10376 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 1492 5899 1544 5908
rect 1492 5865 1501 5899
rect 1501 5865 1535 5899
rect 1535 5865 1544 5899
rect 1492 5856 1544 5865
rect 4160 5856 4212 5908
rect 4804 5856 4856 5908
rect 5540 5856 5592 5908
rect 5632 5856 5684 5908
rect 3700 5788 3752 5840
rect 5264 5788 5316 5840
rect 4160 5720 4212 5772
rect 2596 5695 2648 5704
rect 2596 5661 2625 5695
rect 2625 5661 2648 5695
rect 2596 5652 2648 5661
rect 4436 5652 4488 5704
rect 5724 5788 5776 5840
rect 3516 5584 3568 5636
rect 2688 5516 2740 5568
rect 4436 5516 4488 5568
rect 4712 5584 4764 5636
rect 5724 5652 5776 5704
rect 7380 5899 7432 5908
rect 7380 5865 7389 5899
rect 7389 5865 7423 5899
rect 7423 5865 7432 5899
rect 7380 5856 7432 5865
rect 6184 5720 6236 5772
rect 7104 5788 7156 5840
rect 8944 5788 8996 5840
rect 10048 5856 10100 5908
rect 9404 5831 9456 5840
rect 9404 5797 9413 5831
rect 9413 5797 9447 5831
rect 9447 5797 9456 5831
rect 9404 5788 9456 5797
rect 10232 5788 10284 5840
rect 6552 5720 6604 5772
rect 6276 5584 6328 5636
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7012 5652 7064 5704
rect 9036 5720 9088 5772
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 8852 5652 8904 5704
rect 9220 5652 9272 5704
rect 9864 5652 9916 5704
rect 5724 5559 5776 5568
rect 5724 5525 5733 5559
rect 5733 5525 5767 5559
rect 5767 5525 5776 5559
rect 5724 5516 5776 5525
rect 5816 5516 5868 5568
rect 6092 5559 6144 5568
rect 6092 5525 6117 5559
rect 6117 5525 6144 5559
rect 6092 5516 6144 5525
rect 6460 5559 6512 5568
rect 6460 5525 6469 5559
rect 6469 5525 6503 5559
rect 6503 5525 6512 5559
rect 6460 5516 6512 5525
rect 6736 5516 6788 5568
rect 7380 5584 7432 5636
rect 7656 5584 7708 5636
rect 7748 5584 7800 5636
rect 8024 5584 8076 5636
rect 8392 5584 8444 5636
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 6920 5516 6972 5525
rect 7104 5516 7156 5568
rect 8576 5516 8628 5568
rect 8668 5516 8720 5568
rect 9220 5559 9272 5568
rect 9220 5525 9229 5559
rect 9229 5525 9263 5559
rect 9263 5525 9272 5559
rect 9220 5516 9272 5525
rect 9496 5516 9548 5568
rect 9864 5516 9916 5568
rect 10416 5559 10468 5568
rect 10416 5525 10425 5559
rect 10425 5525 10459 5559
rect 10459 5525 10468 5559
rect 10416 5516 10468 5525
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 1952 5355 2004 5364
rect 1952 5321 1961 5355
rect 1961 5321 1995 5355
rect 1995 5321 2004 5355
rect 1952 5312 2004 5321
rect 5448 5312 5500 5364
rect 5540 5355 5592 5364
rect 5540 5321 5549 5355
rect 5549 5321 5583 5355
rect 5583 5321 5592 5355
rect 5540 5312 5592 5321
rect 5632 5312 5684 5364
rect 6000 5312 6052 5364
rect 1492 5176 1544 5228
rect 2228 5176 2280 5228
rect 4068 5244 4120 5296
rect 3148 5176 3200 5228
rect 4896 5219 4948 5228
rect 4896 5185 4914 5219
rect 4914 5185 4948 5219
rect 4896 5176 4948 5185
rect 2964 5108 3016 5160
rect 3056 5151 3108 5160
rect 3056 5117 3065 5151
rect 3065 5117 3099 5151
rect 3099 5117 3108 5151
rect 3056 5108 3108 5117
rect 5264 5108 5316 5160
rect 6460 5244 6512 5296
rect 6920 5244 6972 5296
rect 7472 5244 7524 5296
rect 6552 5176 6604 5228
rect 5908 5108 5960 5160
rect 1584 4972 1636 5024
rect 2872 4972 2924 5024
rect 3240 4972 3292 5024
rect 4068 4972 4120 5024
rect 5448 5040 5500 5092
rect 5540 5040 5592 5092
rect 6920 5040 6972 5092
rect 6276 4972 6328 5024
rect 6460 4972 6512 5024
rect 7288 4972 7340 5024
rect 8208 5219 8260 5228
rect 8208 5185 8217 5219
rect 8217 5185 8251 5219
rect 8251 5185 8260 5219
rect 8208 5176 8260 5185
rect 9404 5219 9456 5228
rect 10324 5287 10376 5296
rect 10324 5253 10333 5287
rect 10333 5253 10367 5287
rect 10367 5253 10376 5287
rect 10324 5244 10376 5253
rect 9404 5185 9422 5219
rect 9422 5185 9456 5219
rect 9404 5176 9456 5185
rect 8668 5108 8720 5160
rect 8208 4972 8260 5024
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 8300 4972 8352 4981
rect 9956 5015 10008 5024
rect 9956 4981 9965 5015
rect 9965 4981 9999 5015
rect 9999 4981 10008 5015
rect 9956 4972 10008 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 2872 4811 2924 4820
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 4160 4768 4212 4820
rect 4252 4768 4304 4820
rect 3792 4700 3844 4752
rect 5172 4768 5224 4820
rect 7380 4768 7432 4820
rect 8024 4811 8076 4820
rect 8024 4777 8033 4811
rect 8033 4777 8067 4811
rect 8067 4777 8076 4811
rect 8024 4768 8076 4777
rect 8300 4768 8352 4820
rect 10508 4768 10560 4820
rect 3516 4675 3568 4684
rect 3516 4641 3525 4675
rect 3525 4641 3559 4675
rect 3559 4641 3568 4675
rect 3516 4632 3568 4641
rect 3976 4564 4028 4616
rect 4068 4564 4120 4616
rect 3424 4496 3476 4548
rect 4896 4539 4948 4548
rect 3148 4471 3200 4480
rect 3148 4437 3157 4471
rect 3157 4437 3191 4471
rect 3191 4437 3200 4471
rect 3148 4428 3200 4437
rect 4436 4428 4488 4480
rect 4896 4505 4905 4539
rect 4905 4505 4939 4539
rect 4939 4505 4948 4539
rect 4896 4496 4948 4505
rect 5080 4539 5132 4548
rect 5080 4505 5105 4539
rect 5105 4505 5132 4539
rect 5080 4496 5132 4505
rect 5356 4564 5408 4616
rect 6460 4496 6512 4548
rect 9864 4632 9916 4684
rect 7288 4564 7340 4616
rect 6920 4539 6972 4548
rect 6552 4471 6604 4480
rect 6552 4437 6561 4471
rect 6561 4437 6595 4471
rect 6595 4437 6604 4471
rect 6552 4428 6604 4437
rect 6920 4505 6932 4539
rect 6932 4505 6972 4539
rect 6920 4496 6972 4505
rect 7012 4496 7064 4548
rect 9864 4496 9916 4548
rect 10416 4471 10468 4480
rect 10416 4437 10425 4471
rect 10425 4437 10459 4471
rect 10459 4437 10468 4471
rect 10416 4428 10468 4437
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 1492 4224 1544 4276
rect 1216 4088 1268 4140
rect 3148 4224 3200 4276
rect 6000 4224 6052 4276
rect 6552 4224 6604 4276
rect 9680 4224 9732 4276
rect 2412 4199 2464 4208
rect 2412 4165 2421 4199
rect 2421 4165 2455 4199
rect 2455 4165 2464 4199
rect 2412 4156 2464 4165
rect 3056 4156 3108 4208
rect 6092 4156 6144 4208
rect 1400 4020 1452 4072
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 2504 4088 2556 4140
rect 2964 4088 3016 4140
rect 1860 4020 1912 4072
rect 1768 3952 1820 4004
rect 2596 4020 2648 4072
rect 3332 4020 3384 4072
rect 4528 4020 4580 4072
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 5540 4088 5592 4140
rect 6184 4088 6236 4140
rect 5080 4063 5132 4072
rect 5080 4029 5089 4063
rect 5089 4029 5123 4063
rect 5123 4029 5132 4063
rect 5080 4020 5132 4029
rect 4620 3952 4672 4004
rect 4712 3952 4764 4004
rect 5356 4020 5408 4072
rect 6460 4020 6512 4072
rect 6644 4156 6696 4208
rect 6828 4199 6880 4208
rect 6828 4165 6837 4199
rect 6837 4165 6871 4199
rect 6871 4165 6880 4199
rect 6828 4156 6880 4165
rect 7840 4199 7892 4208
rect 7840 4165 7849 4199
rect 7849 4165 7883 4199
rect 7883 4165 7892 4199
rect 7840 4156 7892 4165
rect 8576 4156 8628 4208
rect 1584 3884 1636 3936
rect 2136 3884 2188 3936
rect 2596 3884 2648 3936
rect 2688 3884 2740 3936
rect 3792 3884 3844 3936
rect 5816 3952 5868 4004
rect 5908 3884 5960 3936
rect 7380 3952 7432 4004
rect 8944 3884 8996 3936
rect 10048 3884 10100 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 4804 3723 4856 3732
rect 4804 3689 4813 3723
rect 4813 3689 4847 3723
rect 4847 3689 4856 3723
rect 4804 3680 4856 3689
rect 2044 3587 2096 3596
rect 2044 3553 2053 3587
rect 2053 3553 2087 3587
rect 2087 3553 2096 3587
rect 2044 3544 2096 3553
rect 3608 3544 3660 3596
rect 5264 3544 5316 3596
rect 8484 3680 8536 3732
rect 7196 3655 7248 3664
rect 7196 3621 7205 3655
rect 7205 3621 7239 3655
rect 7239 3621 7248 3655
rect 7196 3612 7248 3621
rect 7380 3655 7432 3664
rect 7380 3621 7389 3655
rect 7389 3621 7423 3655
rect 7423 3621 7432 3655
rect 7380 3612 7432 3621
rect 8300 3612 8352 3664
rect 8116 3544 8168 3596
rect 9772 3680 9824 3732
rect 9864 3723 9916 3732
rect 9864 3689 9873 3723
rect 9873 3689 9907 3723
rect 9907 3689 9916 3723
rect 9864 3680 9916 3689
rect 2412 3408 2464 3460
rect 2688 3408 2740 3460
rect 4896 3476 4948 3528
rect 5448 3476 5500 3528
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 5724 3476 5776 3528
rect 6184 3476 6236 3528
rect 9496 3519 9548 3528
rect 9496 3485 9505 3519
rect 9505 3485 9539 3519
rect 9539 3485 9548 3519
rect 9496 3476 9548 3485
rect 9772 3476 9824 3528
rect 10140 3476 10192 3528
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 10784 3476 10836 3528
rect 6368 3408 6420 3460
rect 6460 3408 6512 3460
rect 6276 3340 6328 3392
rect 6644 3340 6696 3392
rect 9220 3340 9272 3392
rect 10048 3340 10100 3392
rect 10692 3408 10744 3460
rect 10416 3383 10468 3392
rect 10416 3349 10425 3383
rect 10425 3349 10459 3383
rect 10459 3349 10468 3383
rect 10416 3340 10468 3349
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 4160 3136 4212 3188
rect 4988 3136 5040 3188
rect 5816 3136 5868 3188
rect 6736 3136 6788 3188
rect 1676 3043 1728 3052
rect 1676 3009 1710 3043
rect 1710 3009 1728 3043
rect 1676 3000 1728 3009
rect 2504 2932 2556 2984
rect 2964 3000 3016 3052
rect 3148 3000 3200 3052
rect 3792 3000 3844 3052
rect 3976 3000 4028 3052
rect 4712 3068 4764 3120
rect 5080 3068 5132 3120
rect 4160 2796 4212 2848
rect 4896 3000 4948 3052
rect 5632 3000 5684 3052
rect 6276 3000 6328 3052
rect 7288 3136 7340 3188
rect 9036 3136 9088 3188
rect 9220 3136 9272 3188
rect 9404 3179 9456 3188
rect 9404 3145 9413 3179
rect 9413 3145 9447 3179
rect 9447 3145 9456 3179
rect 9404 3136 9456 3145
rect 10876 3068 10928 3120
rect 9128 3000 9180 3052
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 10048 3043 10100 3052
rect 10048 3009 10057 3043
rect 10057 3009 10091 3043
rect 10091 3009 10100 3043
rect 10048 3000 10100 3009
rect 10140 3043 10192 3052
rect 10140 3009 10149 3043
rect 10149 3009 10183 3043
rect 10183 3009 10192 3043
rect 10140 3000 10192 3009
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 5356 2864 5408 2916
rect 10232 2932 10284 2984
rect 5724 2796 5776 2848
rect 6644 2864 6696 2916
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 940 2592 992 2644
rect 756 2456 808 2508
rect 1860 2456 1912 2508
rect 2596 2456 2648 2508
rect 6736 2592 6788 2644
rect 6828 2592 6880 2644
rect 4436 2524 4488 2576
rect 5632 2524 5684 2576
rect 1768 2320 1820 2372
rect 2320 2388 2372 2440
rect 2412 2320 2464 2372
rect 4160 2320 4212 2372
rect 7380 2388 7432 2440
rect 8116 2388 8168 2440
rect 8208 2388 8260 2440
rect 9956 2431 10008 2440
rect 9956 2397 9965 2431
rect 9965 2397 9999 2431
rect 9999 2397 10008 2431
rect 9956 2388 10008 2397
rect 10232 2431 10284 2440
rect 10232 2397 10241 2431
rect 10241 2397 10275 2431
rect 10275 2397 10284 2431
rect 10232 2388 10284 2397
rect 10140 2295 10192 2304
rect 10140 2261 10149 2295
rect 10149 2261 10183 2295
rect 10183 2261 10192 2295
rect 10140 2252 10192 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
rect 10876 2184 10928 2236
rect 756 2048 808 2100
rect 7288 2048 7340 2100
<< metal2 >>
rect 8482 12880 8538 12889
rect 8482 12815 8538 12824
rect 1676 11620 1728 11626
rect 1676 11562 1728 11568
rect 1688 11354 1716 11562
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1768 11280 1820 11286
rect 1490 11248 1546 11257
rect 1768 11222 1820 11228
rect 1490 11183 1546 11192
rect 1584 11212 1636 11218
rect 1504 11150 1532 11183
rect 1584 11154 1636 11160
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 940 9988 992 9994
rect 940 9930 992 9936
rect 664 9580 716 9586
rect 664 9522 716 9528
rect 676 2088 704 9522
rect 756 7200 808 7206
rect 756 7142 808 7148
rect 768 2514 796 7142
rect 952 2650 980 9930
rect 1504 9674 1532 10610
rect 1412 9646 1532 9674
rect 1216 9104 1268 9110
rect 1216 9046 1268 9052
rect 1124 8424 1176 8430
rect 1124 8366 1176 8372
rect 1030 5672 1086 5681
rect 1030 5607 1086 5616
rect 940 2644 992 2650
rect 940 2586 992 2592
rect 756 2508 808 2514
rect 756 2450 808 2456
rect 1044 2281 1072 5607
rect 1136 4049 1164 8366
rect 1228 4146 1256 9046
rect 1308 7948 1360 7954
rect 1308 7890 1360 7896
rect 1320 6712 1348 7890
rect 1412 6780 1440 9646
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1504 6905 1532 7346
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 1412 6752 1532 6780
rect 1320 6684 1440 6712
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1320 4729 1348 6258
rect 1306 4720 1362 4729
rect 1306 4655 1362 4664
rect 1216 4140 1268 4146
rect 1216 4082 1268 4088
rect 1412 4078 1440 6684
rect 1504 6458 1532 6752
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 1492 6180 1544 6186
rect 1492 6122 1544 6128
rect 1504 5914 1532 6122
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1504 4282 1532 5170
rect 1596 5030 1624 11154
rect 1780 10962 1808 11222
rect 2608 11218 2636 11494
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1688 10934 1808 10962
rect 1688 10674 1716 10934
rect 1872 10810 1900 11086
rect 3068 11082 3096 11222
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1674 10568 1730 10577
rect 1674 10503 1730 10512
rect 1688 10062 1716 10503
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1492 4276 1544 4282
rect 1492 4218 1544 4224
rect 1400 4072 1452 4078
rect 1122 4040 1178 4049
rect 1400 4014 1452 4020
rect 1122 3975 1178 3984
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1596 2774 1624 3878
rect 1688 3058 1716 9862
rect 1780 4010 1808 10746
rect 2516 10606 2544 11018
rect 2610 10908 2918 10917
rect 2610 10906 2616 10908
rect 2672 10906 2696 10908
rect 2752 10906 2776 10908
rect 2832 10906 2856 10908
rect 2912 10906 2918 10908
rect 2672 10854 2674 10906
rect 2854 10854 2856 10906
rect 2610 10852 2616 10854
rect 2672 10852 2696 10854
rect 2752 10852 2776 10854
rect 2832 10852 2856 10854
rect 2912 10852 2918 10854
rect 2610 10843 2918 10852
rect 3160 10810 3188 11222
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 1872 9625 1900 10406
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 2332 10033 2360 10406
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2318 10024 2374 10033
rect 2318 9959 2374 9968
rect 2884 9926 2912 10202
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 1858 9616 1914 9625
rect 1858 9551 1914 9560
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2332 9489 2360 9522
rect 2318 9480 2374 9489
rect 2318 9415 2374 9424
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 2320 8900 2372 8906
rect 2320 8842 2372 8848
rect 1950 8392 2006 8401
rect 1872 8350 1950 8378
rect 1872 6458 1900 8350
rect 1950 8327 2006 8336
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2228 6928 2280 6934
rect 1950 6896 2006 6905
rect 2228 6870 2280 6876
rect 1950 6831 2006 6840
rect 1964 6798 1992 6831
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1964 6202 1992 6598
rect 1872 6174 1992 6202
rect 2148 6202 2176 6598
rect 2240 6458 2268 6870
rect 2332 6746 2360 8842
rect 2410 8528 2466 8537
rect 2410 8463 2466 8472
rect 2424 7290 2452 8463
rect 2516 7546 2544 9862
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 2976 9466 3004 9998
rect 2884 9438 3004 9466
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 8945 2820 9318
rect 2884 9042 2912 9438
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2778 8936 2834 8945
rect 2778 8871 2834 8880
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2976 7750 3004 9318
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2424 7262 2636 7290
rect 2502 7168 2558 7177
rect 2502 7103 2558 7112
rect 2516 6866 2544 7103
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2332 6718 2452 6746
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2226 6216 2282 6225
rect 2148 6174 2226 6202
rect 1872 4185 1900 6174
rect 2226 6151 2282 6160
rect 2240 6118 2268 6151
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2226 5808 2282 5817
rect 2226 5743 2282 5752
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1964 5273 1992 5306
rect 1950 5264 2006 5273
rect 2240 5234 2268 5743
rect 1950 5199 2006 5208
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1858 4176 1914 4185
rect 1858 4111 1914 4120
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1768 4004 1820 4010
rect 1768 3946 1820 3952
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1596 2746 1808 2774
rect 1780 2378 1808 2746
rect 1872 2514 1900 4014
rect 2148 3942 2176 4082
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2042 3632 2098 3641
rect 2042 3567 2044 3576
rect 2096 3567 2098 3576
rect 2044 3538 2096 3544
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 2332 2446 2360 6598
rect 2424 6338 2452 6718
rect 2608 6662 2636 7262
rect 2700 7002 2728 7346
rect 2976 7324 3004 7686
rect 3068 7478 3096 10610
rect 3160 10305 3188 10746
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 3146 10296 3202 10305
rect 3146 10231 3202 10240
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3160 8430 3188 9998
rect 3252 9926 3280 10610
rect 3436 10062 3464 11290
rect 3700 11280 3752 11286
rect 3700 11222 3752 11228
rect 3712 11082 3740 11222
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 3700 11076 3752 11082
rect 3700 11018 3752 11024
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3528 10713 3556 10950
rect 3514 10704 3570 10713
rect 3514 10639 3570 10648
rect 3804 10606 3832 11018
rect 3974 10840 4030 10849
rect 3974 10775 4030 10784
rect 4068 10804 4120 10810
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3252 9761 3280 9862
rect 3238 9752 3294 9761
rect 3238 9687 3294 9696
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3160 7721 3188 8366
rect 3146 7712 3202 7721
rect 3146 7647 3202 7656
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 2870 7304 2926 7313
rect 2976 7296 3096 7324
rect 2870 7239 2926 7248
rect 2884 7154 2912 7239
rect 2884 7126 3004 7154
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2870 6896 2926 6905
rect 2870 6831 2926 6840
rect 2688 6792 2740 6798
rect 2686 6760 2688 6769
rect 2740 6760 2742 6769
rect 2686 6695 2742 6704
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2780 6656 2832 6662
rect 2884 6644 2912 6831
rect 2832 6616 2912 6644
rect 2780 6598 2832 6604
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2688 6384 2740 6390
rect 2686 6352 2688 6361
rect 2872 6384 2924 6390
rect 2740 6352 2742 6361
rect 2424 6310 2544 6338
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 4214 2452 6054
rect 2516 4264 2544 6310
rect 2976 6372 3004 7126
rect 2924 6344 3004 6372
rect 2872 6326 2924 6332
rect 2686 6287 2742 6296
rect 2594 5808 2650 5817
rect 2594 5743 2650 5752
rect 2608 5710 2636 5743
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2700 5574 2728 6287
rect 3068 6236 3096 7296
rect 3252 6984 3280 8978
rect 2976 6208 3096 6236
rect 3160 6956 3280 6984
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2976 5166 3004 6208
rect 3160 5953 3188 6956
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3252 6730 3280 6802
rect 3344 6798 3372 9862
rect 3436 9042 3464 9998
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3436 8634 3464 8842
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3436 6905 3464 7686
rect 3422 6896 3478 6905
rect 3422 6831 3478 6840
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3146 5944 3202 5953
rect 3146 5879 3202 5888
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 2964 5160 3016 5166
rect 3056 5160 3108 5166
rect 2964 5102 3016 5108
rect 3054 5128 3056 5137
rect 3108 5128 3110 5137
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2884 4826 2912 4966
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2516 4236 2728 4264
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2424 2378 2452 3402
rect 2516 2990 2544 4082
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2608 3942 2636 4014
rect 2700 3942 2728 4236
rect 2976 4146 3004 5102
rect 3054 5063 3110 5072
rect 3160 5001 3188 5170
rect 3252 5030 3280 6666
rect 3344 5545 3372 6734
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6322 3464 6598
rect 3528 6322 3556 10406
rect 3606 10296 3662 10305
rect 3606 10231 3662 10240
rect 3620 10130 3648 10231
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3712 10062 3740 10406
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3606 9072 3662 9081
rect 3606 9007 3662 9016
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3330 5536 3386 5545
rect 3330 5471 3386 5480
rect 3330 5400 3386 5409
rect 3330 5335 3386 5344
rect 3240 5024 3292 5030
rect 3146 4992 3202 5001
rect 3068 4950 3146 4978
rect 3068 4214 3096 4950
rect 3240 4966 3292 4972
rect 3146 4927 3202 4936
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3160 4282 3188 4422
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3056 4208 3108 4214
rect 3056 4150 3108 4156
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2700 3466 2728 3878
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 3252 3074 3280 4966
rect 3344 4078 3372 5335
rect 3436 4554 3464 6258
rect 3528 6089 3556 6258
rect 3514 6080 3570 6089
rect 3514 6015 3570 6024
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3528 4690 3556 5578
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3424 4548 3476 4554
rect 3424 4490 3476 4496
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3620 3602 3648 9007
rect 3712 7750 3740 9454
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3698 7576 3754 7585
rect 3698 7511 3700 7520
rect 3752 7511 3754 7520
rect 3700 7482 3752 7488
rect 3698 7440 3754 7449
rect 3698 7375 3754 7384
rect 3712 6662 3740 7375
rect 3804 7002 3832 10542
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3896 6866 3924 10610
rect 3988 10266 4016 10775
rect 4068 10746 4120 10752
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3988 9382 4016 10202
rect 4080 10062 4108 10746
rect 4172 10742 4200 11154
rect 4540 11014 4568 11494
rect 6950 11452 7258 11461
rect 6950 11450 6956 11452
rect 7012 11450 7036 11452
rect 7092 11450 7116 11452
rect 7172 11450 7196 11452
rect 7252 11450 7258 11452
rect 7012 11398 7014 11450
rect 7194 11398 7196 11450
rect 6950 11396 6956 11398
rect 7012 11396 7036 11398
rect 7092 11396 7116 11398
rect 7172 11396 7196 11398
rect 7252 11396 7258 11398
rect 6950 11387 7258 11396
rect 8496 11354 8524 12815
rect 9586 11792 9642 11801
rect 9586 11727 9642 11736
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 5644 11132 5672 11222
rect 5724 11144 5776 11150
rect 5644 11121 5724 11132
rect 5630 11112 5724 11121
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 5540 11076 5592 11082
rect 5686 11104 5724 11112
rect 5724 11086 5776 11092
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5630 11047 5686 11056
rect 5540 11018 5592 11024
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4632 10742 4660 11018
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4080 9518 4108 9998
rect 4252 9920 4304 9926
rect 4436 9920 4488 9926
rect 4252 9862 4304 9868
rect 4434 9888 4436 9897
rect 4488 9888 4490 9897
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3988 8809 4016 9318
rect 3974 8800 4030 8809
rect 3974 8735 4030 8744
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3988 8265 4016 8570
rect 4080 8430 4108 9318
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3974 8256 4030 8265
rect 3974 8191 4030 8200
rect 3974 7984 4030 7993
rect 3974 7919 4030 7928
rect 3988 7546 4016 7919
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 4080 7342 4108 8366
rect 4172 8362 4200 9386
rect 4264 8634 4292 9862
rect 4434 9823 4490 9832
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4356 8430 4384 8774
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4342 8256 4398 8265
rect 4342 8191 4398 8200
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4068 7336 4120 7342
rect 3988 7296 4068 7324
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3988 6254 4016 7296
rect 4068 7278 4120 7284
rect 4066 6896 4122 6905
rect 4066 6831 4122 6840
rect 3792 6248 3844 6254
rect 3712 6208 3792 6236
rect 3712 5846 3740 6208
rect 3792 6190 3844 6196
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3700 5840 3752 5846
rect 3700 5782 3752 5788
rect 3804 4758 3832 6054
rect 3896 4865 3924 6054
rect 3974 5944 4030 5953
rect 3974 5879 4030 5888
rect 3882 4856 3938 4865
rect 3882 4791 3938 4800
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3988 4622 4016 5879
rect 4080 5302 4108 6831
rect 4172 5914 4200 7346
rect 4356 6390 4384 8191
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4622 4108 4966
rect 4172 4826 4200 5714
rect 4264 4826 4292 6190
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4356 4298 4384 6326
rect 4448 5710 4476 9522
rect 4540 8537 4568 10202
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4632 9654 4660 9998
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4724 9722 4752 9930
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4620 9648 4672 9654
rect 4672 9596 4752 9602
rect 4620 9590 4752 9596
rect 4632 9574 4752 9590
rect 4724 8566 4752 9574
rect 4816 9110 4844 9998
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4908 9654 4936 9862
rect 5552 9761 5580 11018
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5538 9752 5594 9761
rect 5538 9687 5594 9696
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 5080 9580 5132 9586
rect 5000 9540 5080 9568
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4896 8900 4948 8906
rect 5000 8888 5028 9540
rect 5080 9522 5132 9528
rect 4948 8860 5028 8888
rect 5080 8900 5132 8906
rect 4896 8842 4948 8848
rect 5080 8842 5132 8848
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 4712 8560 4764 8566
rect 4526 8528 4582 8537
rect 4712 8502 4764 8508
rect 4526 8463 4582 8472
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4448 4486 4476 5510
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4356 4270 4476 4298
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 3160 3058 3280 3074
rect 3804 3058 3832 3878
rect 4158 3496 4214 3505
rect 4158 3431 4214 3440
rect 4172 3194 4200 3431
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 3148 3052 3280 3058
rect 3200 3046 3280 3052
rect 3792 3052 3844 3058
rect 3148 2994 3200 3000
rect 3792 2994 3844 3000
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 2504 2984 2556 2990
rect 2976 2961 3004 2994
rect 2504 2926 2556 2932
rect 2962 2952 3018 2961
rect 2516 2774 2544 2926
rect 3988 2938 4016 2994
rect 4066 2952 4122 2961
rect 3988 2910 4066 2938
rect 2962 2887 3018 2896
rect 4066 2887 4122 2896
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 2516 2746 2636 2774
rect 2608 2514 2636 2746
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 4172 2378 4200 2790
rect 4448 2582 4476 4270
rect 4540 4078 4568 8298
rect 4620 7200 4672 7206
rect 4724 7177 4752 8502
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4620 7142 4672 7148
rect 4710 7168 4766 7177
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4632 4010 4660 7142
rect 4710 7103 4766 7112
rect 4724 5642 4752 7103
rect 4816 5914 4844 8230
rect 4908 8090 4936 8842
rect 4896 8084 4948 8090
rect 4948 8044 5028 8072
rect 4896 8026 4948 8032
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4908 6633 4936 7754
rect 4894 6624 4950 6633
rect 4894 6559 4950 6568
rect 4894 6352 4950 6361
rect 4894 6287 4950 6296
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4908 5794 4936 6287
rect 5000 6118 5028 8044
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4816 5766 4936 5794
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4710 5400 4766 5409
rect 4710 5335 4766 5344
rect 4724 4010 4752 5335
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4816 3738 4844 5766
rect 5092 5250 5120 8842
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 4908 5234 5120 5250
rect 4896 5228 5120 5234
rect 4948 5222 5120 5228
rect 4896 5170 4948 5176
rect 5184 4826 5212 8434
rect 5262 8120 5318 8129
rect 5262 8055 5264 8064
rect 5316 8055 5318 8064
rect 5264 8026 5316 8032
rect 5368 7886 5396 8774
rect 5552 8401 5580 8842
rect 5538 8392 5594 8401
rect 5538 8327 5594 8336
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5276 6798 5304 7822
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5276 5846 5304 6734
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5276 5166 5304 5782
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5170 4584 5226 4593
rect 5092 4554 5170 4570
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 5080 4548 5170 4554
rect 5132 4542 5170 4548
rect 5170 4519 5226 4528
rect 5080 4490 5132 4496
rect 4908 4457 4936 4490
rect 4894 4448 4950 4457
rect 4894 4383 4950 4392
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4710 3360 4766 3369
rect 4710 3295 4766 3304
rect 4724 3126 4752 3295
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4908 3058 4936 3470
rect 5000 3194 5028 4082
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5092 3126 5120 4014
rect 5276 3602 5304 5102
rect 5368 4622 5396 7686
rect 5460 7546 5488 8230
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5552 7478 5580 8230
rect 5644 7750 5672 10678
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5460 5681 5488 6666
rect 5552 6390 5580 6938
rect 5644 6458 5672 7686
rect 5736 6798 5764 10950
rect 5828 10674 5856 11086
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7208 10810 7236 10950
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7286 10704 7342 10713
rect 5816 10668 5868 10674
rect 7286 10639 7342 10648
rect 5816 10610 5868 10616
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 6368 10532 6420 10538
rect 6368 10474 6420 10480
rect 6012 9722 6040 10474
rect 6276 10192 6328 10198
rect 6182 10160 6238 10169
rect 6104 10130 6182 10146
rect 6092 10124 6182 10130
rect 6144 10118 6182 10124
rect 6276 10134 6328 10140
rect 6182 10095 6238 10104
rect 6092 10066 6144 10072
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 9042 5856 9318
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5722 6488 5778 6497
rect 5632 6452 5684 6458
rect 5722 6423 5778 6432
rect 5632 6394 5684 6400
rect 5540 6384 5592 6390
rect 5736 6338 5764 6423
rect 5540 6326 5592 6332
rect 5644 6310 5764 6338
rect 5644 6118 5672 6310
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5644 5914 5672 6054
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5446 5672 5502 5681
rect 5446 5607 5502 5616
rect 5552 5370 5580 5850
rect 5736 5846 5764 6054
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5724 5704 5776 5710
rect 5722 5672 5724 5681
rect 5776 5672 5778 5681
rect 5722 5607 5778 5616
rect 5828 5574 5856 8978
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5920 8634 5948 8910
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 6012 8498 6040 9386
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6012 7426 6040 8434
rect 6104 7818 6132 9862
rect 6196 7886 6224 9998
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6092 7812 6144 7818
rect 6092 7754 6144 7760
rect 6012 7398 6224 7426
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 5908 7200 5960 7206
rect 5906 7168 5908 7177
rect 5960 7168 5962 7177
rect 5906 7103 5962 7112
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5724 5568 5776 5574
rect 5630 5536 5686 5545
rect 5724 5510 5776 5516
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5630 5471 5686 5480
rect 5644 5370 5672 5471
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5460 5250 5488 5306
rect 5460 5222 5672 5250
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5354 4312 5410 4321
rect 5354 4247 5410 4256
rect 5368 4078 5396 4247
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 5368 2922 5396 4014
rect 5460 3534 5488 5034
rect 5552 4146 5580 5034
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5538 3768 5594 3777
rect 5538 3703 5594 3712
rect 5552 3534 5580 3703
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5644 3058 5672 5222
rect 5736 3534 5764 5510
rect 5814 5400 5870 5409
rect 5814 5335 5870 5344
rect 5828 4010 5856 5335
rect 5920 5166 5948 6802
rect 6012 5370 6040 7278
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6104 6390 6132 6734
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 6196 6338 6224 7398
rect 6288 6905 6316 10134
rect 6274 6896 6330 6905
rect 6380 6866 6408 10474
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6472 8786 6500 10406
rect 6950 10364 7258 10373
rect 6950 10362 6956 10364
rect 7012 10362 7036 10364
rect 7092 10362 7116 10364
rect 7172 10362 7196 10364
rect 7252 10362 7258 10364
rect 7012 10310 7014 10362
rect 7194 10310 7196 10362
rect 6950 10308 6956 10310
rect 7012 10308 7036 10310
rect 7092 10308 7116 10310
rect 7172 10308 7196 10310
rect 7252 10308 7258 10310
rect 6950 10299 7258 10308
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6656 9654 6684 9998
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6656 8974 6684 9590
rect 6932 9586 6960 9930
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6748 8786 6776 8910
rect 6472 8758 6776 8786
rect 6274 6831 6330 6840
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6472 6458 6500 8758
rect 6734 7984 6790 7993
rect 6840 7970 6868 9318
rect 6950 9276 7258 9285
rect 6950 9274 6956 9276
rect 7012 9274 7036 9276
rect 7092 9274 7116 9276
rect 7172 9274 7196 9276
rect 7252 9274 7258 9276
rect 7012 9222 7014 9274
rect 7194 9222 7196 9274
rect 6950 9220 6956 9222
rect 7012 9220 7036 9222
rect 7092 9220 7116 9222
rect 7172 9220 7196 9222
rect 7252 9220 7258 9222
rect 6950 9211 7258 9220
rect 7300 9042 7328 10639
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8362 6960 8774
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6950 8188 7258 8197
rect 6950 8186 6956 8188
rect 7012 8186 7036 8188
rect 7092 8186 7116 8188
rect 7172 8186 7196 8188
rect 7252 8186 7258 8188
rect 7012 8134 7014 8186
rect 7194 8134 7196 8186
rect 6950 8132 6956 8134
rect 7012 8132 7036 8134
rect 7092 8132 7116 8134
rect 7172 8132 7196 8134
rect 7252 8132 7258 8134
rect 6950 8123 7258 8132
rect 6790 7942 6868 7970
rect 7288 7948 7340 7954
rect 6734 7919 6790 7928
rect 7288 7890 7340 7896
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6564 6730 6592 7822
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6656 7274 6684 7754
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6196 6310 6500 6338
rect 6472 6254 6500 6310
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6472 6100 6500 6190
rect 6380 6072 6500 6100
rect 6274 5944 6330 5953
rect 6274 5879 6330 5888
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6196 5522 6224 5714
rect 6288 5642 6316 5879
rect 6276 5636 6328 5642
rect 6276 5578 6328 5584
rect 6274 5536 6330 5545
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 6012 4282 6040 5306
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 6104 4214 6132 5510
rect 6196 5494 6274 5522
rect 6274 5471 6330 5480
rect 6288 5030 6316 5471
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6092 4208 6144 4214
rect 5906 4176 5962 4185
rect 6092 4150 6144 4156
rect 5906 4111 5962 4120
rect 6184 4140 6236 4146
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 5920 3942 5948 4111
rect 6184 4082 6236 4088
rect 5908 3936 5960 3942
rect 5814 3904 5870 3913
rect 5908 3878 5960 3884
rect 5814 3839 5870 3848
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5828 3194 5856 3839
rect 6196 3534 6224 4082
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6380 3466 6408 6072
rect 6564 5778 6592 6666
rect 6656 6458 6684 6802
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6748 6390 6776 7822
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6840 7002 6868 7346
rect 6932 7313 6960 7754
rect 6918 7304 6974 7313
rect 6918 7239 6974 7248
rect 7300 7154 7328 7890
rect 7392 7478 7420 9862
rect 7484 7546 7512 11018
rect 7610 10908 7918 10917
rect 7610 10906 7616 10908
rect 7672 10906 7696 10908
rect 7752 10906 7776 10908
rect 7832 10906 7856 10908
rect 7912 10906 7918 10908
rect 7672 10854 7674 10906
rect 7854 10854 7856 10906
rect 7610 10852 7616 10854
rect 7672 10852 7696 10854
rect 7752 10852 7776 10854
rect 7832 10852 7856 10854
rect 7912 10852 7918 10854
rect 7610 10843 7918 10852
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7668 10130 7696 10610
rect 7852 10266 7880 10610
rect 7944 10266 7972 10746
rect 8404 10674 8432 11222
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 8114 10568 8170 10577
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7944 9908 7972 10202
rect 8036 10062 8064 10542
rect 8114 10503 8170 10512
rect 8208 10532 8260 10538
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 7944 9880 8064 9908
rect 7610 9820 7918 9829
rect 7610 9818 7616 9820
rect 7672 9818 7696 9820
rect 7752 9818 7776 9820
rect 7832 9818 7856 9820
rect 7912 9818 7918 9820
rect 7672 9766 7674 9818
rect 7854 9766 7856 9818
rect 7610 9764 7616 9766
rect 7672 9764 7696 9766
rect 7752 9764 7776 9766
rect 7832 9764 7856 9766
rect 7912 9764 7918 9766
rect 7610 9755 7918 9764
rect 8036 9722 8064 9880
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7576 8945 7604 9658
rect 8128 9586 8156 10503
rect 8208 10474 8260 10480
rect 8220 9738 8248 10474
rect 8312 10130 8340 10610
rect 8496 10538 8524 11086
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 8496 10266 8524 10474
rect 8588 10266 8616 11562
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8772 10713 8800 11222
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9416 10742 9444 11018
rect 9600 10810 9628 11727
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9404 10736 9456 10742
rect 8758 10704 8814 10713
rect 8668 10668 8720 10674
rect 9404 10678 9456 10684
rect 8758 10639 8814 10648
rect 8668 10610 8720 10616
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8312 9926 8340 10066
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8220 9710 8432 9738
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 7668 9178 7696 9522
rect 7838 9480 7894 9489
rect 7838 9415 7840 9424
rect 7892 9415 7894 9424
rect 7840 9386 7892 9392
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 8036 9081 8064 9318
rect 8022 9072 8078 9081
rect 8022 9007 8078 9016
rect 8024 8968 8076 8974
rect 7562 8936 7618 8945
rect 8024 8910 8076 8916
rect 7562 8871 7618 8880
rect 7610 8732 7918 8741
rect 7610 8730 7616 8732
rect 7672 8730 7696 8732
rect 7752 8730 7776 8732
rect 7832 8730 7856 8732
rect 7912 8730 7918 8732
rect 7672 8678 7674 8730
rect 7854 8678 7856 8730
rect 7610 8676 7616 8678
rect 7672 8676 7696 8678
rect 7752 8676 7776 8678
rect 7832 8676 7856 8678
rect 7912 8676 7918 8678
rect 7610 8667 7918 8676
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7564 7200 7616 7206
rect 7300 7126 7512 7154
rect 7564 7142 7616 7148
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7392 6866 7420 6938
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 6826 6624 6882 6633
rect 6826 6559 6882 6568
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6642 6216 6698 6225
rect 6748 6202 6776 6326
rect 6840 6225 6868 6559
rect 6918 6488 6974 6497
rect 6918 6423 6974 6432
rect 6932 6390 6960 6423
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 7104 6248 7156 6254
rect 6698 6174 6776 6202
rect 6826 6216 6882 6225
rect 6642 6151 6698 6160
rect 7104 6190 7156 6196
rect 6826 6151 6882 6160
rect 6642 6080 6698 6089
rect 6642 6015 6698 6024
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6472 5302 6500 5510
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6472 4554 6500 4966
rect 6564 4865 6592 5170
rect 6550 4856 6606 4865
rect 6550 4791 6606 4800
rect 6460 4548 6512 4554
rect 6460 4490 6512 4496
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6564 4282 6592 4422
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6656 4214 6684 6015
rect 6840 5794 6868 6151
rect 7116 6100 7144 6190
rect 7116 6072 7328 6100
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 7104 5840 7156 5846
rect 6840 5766 7052 5794
rect 7104 5782 7156 5788
rect 7024 5710 7052 5766
rect 6920 5704 6972 5710
rect 6840 5652 6920 5658
rect 6840 5646 6972 5652
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6840 5630 6960 5646
rect 6736 5568 6788 5574
rect 6734 5536 6736 5545
rect 6788 5536 6790 5545
rect 6734 5471 6790 5480
rect 6734 4992 6790 5001
rect 6840 4978 6868 5630
rect 7116 5574 7144 5782
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 6932 5302 6960 5510
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6932 5098 6960 5238
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 7300 5030 7328 6072
rect 7392 5914 7420 6802
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 6790 4950 6868 4978
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 6734 4927 6790 4936
rect 6840 4740 6868 4950
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 6840 4712 7052 4740
rect 7024 4554 7052 4712
rect 7300 4622 7328 4966
rect 7392 4826 7420 5578
rect 7484 5302 7512 7126
rect 7576 6905 7604 7142
rect 7562 6896 7618 6905
rect 7562 6831 7618 6840
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7610 6491 7918 6500
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7668 5642 7696 6326
rect 7760 5642 7788 6326
rect 7656 5636 7708 5642
rect 7656 5578 7708 5584
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7944 5522 7972 6394
rect 8036 5642 8064 8910
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 7944 5494 8064 5522
rect 7610 5468 7918 5477
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7610 5403 7918 5412
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 8036 4826 8064 5494
rect 8128 4842 8156 8842
rect 8220 7857 8248 9318
rect 8312 9178 8340 9590
rect 8404 9178 8432 9710
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 8362 8340 8910
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8298 7984 8354 7993
rect 8298 7919 8300 7928
rect 8352 7919 8354 7928
rect 8300 7890 8352 7896
rect 8206 7848 8262 7857
rect 8206 7783 8262 7792
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8220 6798 8248 7482
rect 8312 7410 8340 7754
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8220 6458 8248 6734
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8206 5536 8262 5545
rect 8206 5471 8262 5480
rect 8220 5234 8248 5471
rect 8312 5273 8340 6734
rect 8404 5642 8432 8774
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8496 6254 8524 8570
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8588 6186 8616 9386
rect 8680 7886 8708 10610
rect 9126 10568 9182 10577
rect 9126 10503 9182 10512
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8758 8120 8814 8129
rect 8758 8055 8760 8064
rect 8812 8055 8814 8064
rect 8760 8026 8812 8032
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8668 7880 8720 7886
rect 8772 7857 8800 7890
rect 8668 7822 8720 7828
rect 8758 7848 8814 7857
rect 8680 7002 8708 7822
rect 8758 7783 8814 7792
rect 8760 7744 8812 7750
rect 8758 7712 8760 7721
rect 8812 7712 8814 7721
rect 8758 7647 8814 7656
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8666 6624 8722 6633
rect 8666 6559 8722 6568
rect 8680 6458 8708 6559
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8666 6352 8722 6361
rect 8666 6287 8722 6296
rect 8576 6180 8628 6186
rect 8576 6122 8628 6128
rect 8482 6080 8538 6089
rect 8482 6015 8538 6024
rect 8496 5681 8524 6015
rect 8680 5681 8708 6287
rect 8772 5710 8800 7142
rect 8864 5710 8892 10406
rect 8956 8634 8984 10406
rect 9140 10062 9168 10503
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9048 8294 9076 9998
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9232 9722 9260 9862
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9140 9382 9168 9590
rect 9416 9518 9444 10678
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9220 9444 9272 9450
rect 9220 9386 9272 9392
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9140 8498 9168 9318
rect 9232 9178 9260 9386
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 8956 8266 9076 8294
rect 8956 8090 8984 8266
rect 9232 8265 9260 8910
rect 9416 8294 9444 9454
rect 9600 8974 9628 9862
rect 9692 9568 9720 11290
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9876 9994 9904 10202
rect 9954 10160 10010 10169
rect 9954 10095 10010 10104
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9784 9674 9812 9930
rect 9784 9646 9904 9674
rect 9772 9580 9824 9586
rect 9692 9540 9772 9568
rect 9772 9522 9824 9528
rect 9784 9489 9812 9522
rect 9770 9480 9826 9489
rect 9770 9415 9826 9424
rect 9876 9382 9904 9646
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9496 8832 9548 8838
rect 9692 8786 9720 9318
rect 9496 8774 9548 8780
rect 9404 8288 9456 8294
rect 9218 8256 9274 8265
rect 9404 8230 9456 8236
rect 9218 8191 9274 8200
rect 9310 8120 9366 8129
rect 8944 8084 8996 8090
rect 9310 8055 9366 8064
rect 8944 8026 8996 8032
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8956 7546 8984 7890
rect 9218 7848 9274 7857
rect 9140 7806 9218 7834
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 8956 6730 8984 7210
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8956 6458 8984 6666
rect 9140 6458 9168 7806
rect 9218 7783 9274 7792
rect 9220 7744 9272 7750
rect 9218 7712 9220 7721
rect 9272 7712 9274 7721
rect 9218 7647 9274 7656
rect 9324 7274 9352 8055
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9416 7206 9444 8230
rect 9508 7342 9536 8774
rect 9600 8758 9720 8786
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9404 7200 9456 7206
rect 9600 7154 9628 8758
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9404 7142 9456 7148
rect 9508 7126 9628 7154
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8956 5846 8984 6054
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8760 5704 8812 5710
rect 8482 5672 8538 5681
rect 8392 5636 8444 5642
rect 8482 5607 8538 5616
rect 8666 5672 8722 5681
rect 8760 5646 8812 5652
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8666 5607 8722 5616
rect 8392 5578 8444 5584
rect 8298 5264 8354 5273
rect 8208 5228 8260 5234
rect 8298 5199 8354 5208
rect 8208 5170 8260 5176
rect 8206 5128 8262 5137
rect 8206 5063 8262 5072
rect 8220 5030 8248 5063
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 8024 4820 8076 4826
rect 8128 4814 8248 4842
rect 8312 4826 8340 4966
rect 8024 4762 8076 4768
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 6826 4448 6882 4457
rect 6826 4383 6882 4392
rect 6840 4214 6868 4383
rect 6644 4208 6696 4214
rect 6828 4208 6880 4214
rect 6644 4150 6696 4156
rect 6748 4168 6828 4196
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6472 3466 6500 4014
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5644 2582 5672 2994
rect 5724 2848 5776 2854
rect 5828 2836 5856 3130
rect 6288 3058 6316 3334
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6656 2922 6684 3334
rect 6748 3194 6776 4168
rect 6828 4150 6880 4156
rect 6932 3924 6960 4490
rect 6840 3896 6960 3924
rect 6840 3720 6868 3896
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 6840 3692 6960 3720
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 5776 2808 5856 2836
rect 5724 2790 5776 2796
rect 6748 2650 6776 3130
rect 6932 2938 6960 3692
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7208 3074 7236 3606
rect 7300 3194 7328 4558
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 7840 4208 7892 4214
rect 7838 4176 7840 4185
rect 7892 4176 7894 4185
rect 7838 4111 7894 4120
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7392 3670 7420 3946
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7208 3046 7328 3074
rect 6840 2910 6960 2938
rect 6840 2650 6868 2910
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 6950 2683 7258 2692
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 4436 2576 4488 2582
rect 4436 2518 4488 2524
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 1768 2372 1820 2378
rect 1768 2314 1820 2320
rect 2412 2372 2464 2378
rect 2412 2314 2464 2320
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 1030 2272 1086 2281
rect 1030 2207 1086 2216
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 7300 2106 7328 3046
rect 7392 2446 7420 3606
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 8128 2446 8156 3538
rect 8220 2446 8248 4814
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8312 3670 8340 4762
rect 8496 3738 8524 5607
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8588 4214 8616 5510
rect 8680 5166 8708 5510
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8956 3942 8984 5782
rect 9048 5778 9076 6326
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8300 3664 8352 3670
rect 8300 3606 8352 3612
rect 9048 3194 9076 5714
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9140 3058 9168 6394
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9232 6225 9260 6326
rect 9218 6216 9274 6225
rect 9218 6151 9274 6160
rect 9220 5704 9272 5710
rect 9218 5672 9220 5681
rect 9272 5672 9274 5681
rect 9218 5607 9274 5616
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9232 3641 9260 5510
rect 9324 5114 9352 6734
rect 9404 6248 9456 6254
rect 9402 6216 9404 6225
rect 9456 6216 9458 6225
rect 9402 6151 9458 6160
rect 9508 6118 9536 7126
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9416 5930 9444 6054
rect 9416 5902 9536 5930
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 9416 5234 9444 5782
rect 9508 5574 9536 5902
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9324 5086 9536 5114
rect 9402 4040 9458 4049
rect 9402 3975 9458 3984
rect 9218 3632 9274 3641
rect 9218 3567 9274 3576
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9232 3194 9260 3334
rect 9416 3194 9444 3975
rect 9508 3534 9536 5086
rect 9600 4593 9628 6598
rect 9586 4584 9642 4593
rect 9586 4519 9642 4528
rect 9692 4282 9720 8434
rect 9784 6390 9812 9318
rect 9968 8974 9996 10095
rect 10060 9586 10088 10950
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10324 9648 10376 9654
rect 10138 9616 10194 9625
rect 10048 9580 10100 9586
rect 10324 9590 10376 9596
rect 10138 9551 10194 9560
rect 10048 9522 10100 9528
rect 10152 9382 10180 9551
rect 10140 9376 10192 9382
rect 10046 9344 10102 9353
rect 10140 9318 10192 9324
rect 10046 9279 10102 9288
rect 10060 9178 10088 9279
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 9876 8514 9904 8774
rect 9876 8486 9996 8514
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9784 3738 9812 6326
rect 9876 5710 9904 8298
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9876 4690 9904 5510
rect 9968 5114 9996 8486
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 7002 10088 8230
rect 10152 7449 10180 8774
rect 10138 7440 10194 7449
rect 10138 7375 10194 7384
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10244 6882 10272 8842
rect 10336 7546 10364 9590
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10428 8537 10456 9318
rect 10414 8528 10470 8537
rect 10414 8463 10470 8472
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10428 8129 10456 8230
rect 10414 8120 10470 8129
rect 10414 8055 10470 8064
rect 10414 7984 10470 7993
rect 10414 7919 10470 7928
rect 10428 7886 10456 7919
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10428 7449 10456 7686
rect 10414 7440 10470 7449
rect 10414 7375 10470 7384
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 10336 7177 10364 7210
rect 10322 7168 10378 7177
rect 10322 7103 10378 7112
rect 10060 6854 10272 6882
rect 10322 6896 10378 6905
rect 10060 5914 10088 6854
rect 10322 6831 10378 6840
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9968 5086 10088 5114
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9968 4729 9996 4966
rect 9954 4720 10010 4729
rect 9864 4684 9916 4690
rect 9954 4655 10010 4664
rect 9864 4626 9916 4632
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9876 3738 9904 4490
rect 10060 3942 10088 5086
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 10152 3534 10180 6666
rect 10244 6390 10272 6734
rect 10336 6458 10364 6831
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10232 6384 10284 6390
rect 10428 6361 10456 6598
rect 10232 6326 10284 6332
rect 10414 6352 10470 6361
rect 10414 6287 10470 6296
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10232 5840 10284 5846
rect 10230 5808 10232 5817
rect 10284 5808 10286 5817
rect 10230 5743 10286 5752
rect 10336 5302 10364 6054
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10324 5296 10376 5302
rect 10428 5273 10456 5510
rect 10324 5238 10376 5244
rect 10414 5264 10470 5273
rect 10414 5199 10470 5208
rect 10520 4826 10548 9658
rect 10600 7812 10652 7818
rect 10600 7754 10652 7760
rect 10612 7410 10640 7754
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10428 4185 10456 4422
rect 10414 4176 10470 4185
rect 10414 4111 10470 4120
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9784 3058 9812 3470
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10060 3058 10088 3334
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10060 2774 10088 2994
rect 9968 2746 10088 2774
rect 10152 2774 10180 2994
rect 10244 2990 10272 3470
rect 10704 3466 10732 9862
rect 10796 3534 10824 9862
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10428 3097 10456 3334
rect 10888 3126 10916 10202
rect 10876 3120 10928 3126
rect 10414 3088 10470 3097
rect 10324 3052 10376 3058
rect 10876 3062 10928 3068
rect 10414 3023 10470 3032
rect 10324 2994 10376 3000
rect 10232 2984 10284 2990
rect 10336 2961 10364 2994
rect 10232 2926 10284 2932
rect 10322 2952 10378 2961
rect 10322 2887 10378 2896
rect 10152 2746 10272 2774
rect 9968 2446 9996 2746
rect 10244 2446 10272 2746
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 7610 2204 7918 2213
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 756 2100 808 2106
rect 676 2060 756 2088
rect 756 2042 808 2048
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 10152 2009 10180 2246
rect 10876 2236 10928 2242
rect 10876 2178 10928 2184
rect 10138 2000 10194 2009
rect 10138 1935 10194 1944
rect 10888 921 10916 2178
rect 10874 912 10930 921
rect 10874 847 10930 856
<< via2 >>
rect 8482 12824 8538 12880
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 1490 11192 1546 11248
rect 1030 5616 1086 5672
rect 1490 6840 1546 6896
rect 1306 4664 1362 4720
rect 1674 10512 1730 10568
rect 1122 3984 1178 4040
rect 2616 10906 2672 10908
rect 2696 10906 2752 10908
rect 2776 10906 2832 10908
rect 2856 10906 2912 10908
rect 2616 10854 2662 10906
rect 2662 10854 2672 10906
rect 2696 10854 2726 10906
rect 2726 10854 2738 10906
rect 2738 10854 2752 10906
rect 2776 10854 2790 10906
rect 2790 10854 2802 10906
rect 2802 10854 2832 10906
rect 2856 10854 2866 10906
rect 2866 10854 2912 10906
rect 2616 10852 2672 10854
rect 2696 10852 2752 10854
rect 2776 10852 2832 10854
rect 2856 10852 2912 10854
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 2318 9968 2374 10024
rect 1858 9560 1914 9616
rect 2318 9424 2374 9480
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 1950 8336 2006 8392
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1950 6840 2006 6896
rect 2410 8472 2466 8528
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 2778 8880 2834 8936
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 2502 7112 2558 7168
rect 2226 6160 2282 6216
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2226 5752 2282 5808
rect 1950 5208 2006 5264
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1858 4120 1914 4176
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2042 3596 2098 3632
rect 2042 3576 2044 3596
rect 2044 3576 2096 3596
rect 2096 3576 2098 3596
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 3146 10240 3202 10296
rect 3514 10648 3570 10704
rect 3974 10784 4030 10840
rect 3238 9696 3294 9752
rect 3146 7656 3202 7712
rect 2870 7248 2926 7304
rect 2870 6840 2926 6896
rect 2686 6740 2688 6760
rect 2688 6740 2740 6760
rect 2740 6740 2742 6760
rect 2686 6704 2742 6740
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2686 6332 2688 6352
rect 2688 6332 2740 6352
rect 2740 6332 2742 6352
rect 2686 6296 2742 6332
rect 2594 5752 2650 5808
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 3422 6840 3478 6896
rect 3146 5888 3202 5944
rect 3054 5108 3056 5128
rect 3056 5108 3108 5128
rect 3108 5108 3110 5128
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 3054 5072 3110 5108
rect 3606 10240 3662 10296
rect 3606 9016 3662 9072
rect 3330 5480 3386 5536
rect 3330 5344 3386 5400
rect 3146 4936 3202 4992
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 3514 6024 3570 6080
rect 3698 7540 3754 7576
rect 3698 7520 3700 7540
rect 3700 7520 3752 7540
rect 3752 7520 3754 7540
rect 3698 7384 3754 7440
rect 6956 11450 7012 11452
rect 7036 11450 7092 11452
rect 7116 11450 7172 11452
rect 7196 11450 7252 11452
rect 6956 11398 7002 11450
rect 7002 11398 7012 11450
rect 7036 11398 7066 11450
rect 7066 11398 7078 11450
rect 7078 11398 7092 11450
rect 7116 11398 7130 11450
rect 7130 11398 7142 11450
rect 7142 11398 7172 11450
rect 7196 11398 7206 11450
rect 7206 11398 7252 11450
rect 6956 11396 7012 11398
rect 7036 11396 7092 11398
rect 7116 11396 7172 11398
rect 7196 11396 7252 11398
rect 9586 11736 9642 11792
rect 5630 11056 5686 11112
rect 4434 9868 4436 9888
rect 4436 9868 4488 9888
rect 4488 9868 4490 9888
rect 3974 8744 4030 8800
rect 3974 8200 4030 8256
rect 3974 7928 4030 7984
rect 4434 9832 4490 9868
rect 4342 8200 4398 8256
rect 4066 6840 4122 6896
rect 3974 5888 4030 5944
rect 3882 4800 3938 4856
rect 5538 9696 5594 9752
rect 4526 8472 4582 8528
rect 4158 3440 4214 3496
rect 2962 2896 3018 2952
rect 4066 2896 4122 2952
rect 4710 7112 4766 7168
rect 4894 6568 4950 6624
rect 4894 6296 4950 6352
rect 4710 5344 4766 5400
rect 5262 8084 5318 8120
rect 5262 8064 5264 8084
rect 5264 8064 5316 8084
rect 5316 8064 5318 8084
rect 5538 8336 5594 8392
rect 5170 4528 5226 4584
rect 4894 4392 4950 4448
rect 4710 3304 4766 3360
rect 7286 10648 7342 10704
rect 6182 10104 6238 10160
rect 5722 6432 5778 6488
rect 5446 5616 5502 5672
rect 5722 5652 5724 5672
rect 5724 5652 5776 5672
rect 5776 5652 5778 5672
rect 5722 5616 5778 5652
rect 5906 7148 5908 7168
rect 5908 7148 5960 7168
rect 5960 7148 5962 7168
rect 5906 7112 5962 7148
rect 5630 5480 5686 5536
rect 5354 4256 5410 4312
rect 5538 3712 5594 3768
rect 5814 5344 5870 5400
rect 6274 6840 6330 6896
rect 6956 10362 7012 10364
rect 7036 10362 7092 10364
rect 7116 10362 7172 10364
rect 7196 10362 7252 10364
rect 6956 10310 7002 10362
rect 7002 10310 7012 10362
rect 7036 10310 7066 10362
rect 7066 10310 7078 10362
rect 7078 10310 7092 10362
rect 7116 10310 7130 10362
rect 7130 10310 7142 10362
rect 7142 10310 7172 10362
rect 7196 10310 7206 10362
rect 7206 10310 7252 10362
rect 6956 10308 7012 10310
rect 7036 10308 7092 10310
rect 7116 10308 7172 10310
rect 7196 10308 7252 10310
rect 6734 7928 6790 7984
rect 6956 9274 7012 9276
rect 7036 9274 7092 9276
rect 7116 9274 7172 9276
rect 7196 9274 7252 9276
rect 6956 9222 7002 9274
rect 7002 9222 7012 9274
rect 7036 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7092 9274
rect 7116 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7172 9274
rect 7196 9222 7206 9274
rect 7206 9222 7252 9274
rect 6956 9220 7012 9222
rect 7036 9220 7092 9222
rect 7116 9220 7172 9222
rect 7196 9220 7252 9222
rect 6956 8186 7012 8188
rect 7036 8186 7092 8188
rect 7116 8186 7172 8188
rect 7196 8186 7252 8188
rect 6956 8134 7002 8186
rect 7002 8134 7012 8186
rect 7036 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7092 8186
rect 7116 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7172 8186
rect 7196 8134 7206 8186
rect 7206 8134 7252 8186
rect 6956 8132 7012 8134
rect 7036 8132 7092 8134
rect 7116 8132 7172 8134
rect 7196 8132 7252 8134
rect 6274 5888 6330 5944
rect 6274 5480 6330 5536
rect 5906 4120 5962 4176
rect 5814 3848 5870 3904
rect 6918 7248 6974 7304
rect 7616 10906 7672 10908
rect 7696 10906 7752 10908
rect 7776 10906 7832 10908
rect 7856 10906 7912 10908
rect 7616 10854 7662 10906
rect 7662 10854 7672 10906
rect 7696 10854 7726 10906
rect 7726 10854 7738 10906
rect 7738 10854 7752 10906
rect 7776 10854 7790 10906
rect 7790 10854 7802 10906
rect 7802 10854 7832 10906
rect 7856 10854 7866 10906
rect 7866 10854 7912 10906
rect 7616 10852 7672 10854
rect 7696 10852 7752 10854
rect 7776 10852 7832 10854
rect 7856 10852 7912 10854
rect 8114 10512 8170 10568
rect 7616 9818 7672 9820
rect 7696 9818 7752 9820
rect 7776 9818 7832 9820
rect 7856 9818 7912 9820
rect 7616 9766 7662 9818
rect 7662 9766 7672 9818
rect 7696 9766 7726 9818
rect 7726 9766 7738 9818
rect 7738 9766 7752 9818
rect 7776 9766 7790 9818
rect 7790 9766 7802 9818
rect 7802 9766 7832 9818
rect 7856 9766 7866 9818
rect 7866 9766 7912 9818
rect 7616 9764 7672 9766
rect 7696 9764 7752 9766
rect 7776 9764 7832 9766
rect 7856 9764 7912 9766
rect 8758 10648 8814 10704
rect 7838 9444 7894 9480
rect 7838 9424 7840 9444
rect 7840 9424 7892 9444
rect 7892 9424 7894 9444
rect 8022 9016 8078 9072
rect 7562 8880 7618 8936
rect 7616 8730 7672 8732
rect 7696 8730 7752 8732
rect 7776 8730 7832 8732
rect 7856 8730 7912 8732
rect 7616 8678 7662 8730
rect 7662 8678 7672 8730
rect 7696 8678 7726 8730
rect 7726 8678 7738 8730
rect 7738 8678 7752 8730
rect 7776 8678 7790 8730
rect 7790 8678 7802 8730
rect 7802 8678 7832 8730
rect 7856 8678 7866 8730
rect 7866 8678 7912 8730
rect 7616 8676 7672 8678
rect 7696 8676 7752 8678
rect 7776 8676 7832 8678
rect 7856 8676 7912 8678
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 6826 6568 6882 6624
rect 6642 6160 6698 6216
rect 6918 6432 6974 6488
rect 6826 6160 6882 6216
rect 6642 6024 6698 6080
rect 6550 4800 6606 4856
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 6734 5516 6736 5536
rect 6736 5516 6788 5536
rect 6788 5516 6790 5536
rect 6734 5480 6790 5516
rect 6734 4936 6790 4992
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 7562 6840 7618 6896
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 8298 7948 8354 7984
rect 8298 7928 8300 7948
rect 8300 7928 8352 7948
rect 8352 7928 8354 7948
rect 8206 7792 8262 7848
rect 8206 5480 8262 5536
rect 9126 10512 9182 10568
rect 8758 8084 8814 8120
rect 8758 8064 8760 8084
rect 8760 8064 8812 8084
rect 8812 8064 8814 8084
rect 8758 7792 8814 7848
rect 8758 7692 8760 7712
rect 8760 7692 8812 7712
rect 8812 7692 8814 7712
rect 8758 7656 8814 7692
rect 8666 6568 8722 6624
rect 8666 6296 8722 6352
rect 8482 6024 8538 6080
rect 9954 10104 10010 10160
rect 9770 9424 9826 9480
rect 9218 8200 9274 8256
rect 9310 8064 9366 8120
rect 9218 7792 9274 7848
rect 9218 7692 9220 7712
rect 9220 7692 9272 7712
rect 9272 7692 9274 7712
rect 9218 7656 9274 7692
rect 8482 5616 8538 5672
rect 8666 5616 8722 5672
rect 8298 5208 8354 5264
rect 8206 5072 8262 5128
rect 6826 4392 6882 4448
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 7838 4156 7840 4176
rect 7840 4156 7892 4176
rect 7892 4156 7894 4176
rect 7838 4120 7894 4156
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 1030 2216 1086 2272
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 9218 6160 9274 6216
rect 9218 5652 9220 5672
rect 9220 5652 9272 5672
rect 9272 5652 9274 5672
rect 9218 5616 9274 5652
rect 9402 6196 9404 6216
rect 9404 6196 9456 6216
rect 9456 6196 9458 6216
rect 9402 6160 9458 6196
rect 9402 3984 9458 4040
rect 9218 3576 9274 3632
rect 9586 4528 9642 4584
rect 10138 9560 10194 9616
rect 10046 9288 10102 9344
rect 10138 7384 10194 7440
rect 10414 8472 10470 8528
rect 10414 8064 10470 8120
rect 10414 7928 10470 7984
rect 10414 7384 10470 7440
rect 10322 7112 10378 7168
rect 10322 6840 10378 6896
rect 9954 4664 10010 4720
rect 10414 6296 10470 6352
rect 10230 5788 10232 5808
rect 10232 5788 10284 5808
rect 10284 5788 10286 5808
rect 10230 5752 10286 5788
rect 10414 5208 10470 5264
rect 10414 4120 10470 4176
rect 10414 3032 10470 3088
rect 10322 2896 10378 2952
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
rect 10138 1944 10194 2000
rect 10874 856 10930 912
<< metal3 >>
rect 8477 12882 8543 12885
rect 11108 12882 11908 12912
rect 8477 12880 11908 12882
rect 8477 12824 8482 12880
rect 8538 12824 11908 12880
rect 8477 12822 11908 12824
rect 8477 12819 8543 12822
rect 11108 12792 11908 12822
rect 9581 11794 9647 11797
rect 11108 11794 11908 11824
rect 9581 11792 11908 11794
rect 9581 11736 9586 11792
rect 9642 11736 11908 11792
rect 9581 11734 11908 11736
rect 9581 11731 9647 11734
rect 11108 11704 11908 11734
rect 0 11524 800 11552
rect 0 11460 796 11524
rect 860 11460 866 11524
rect 0 11432 800 11460
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 6946 11456 7262 11457
rect 6946 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7262 11456
rect 6946 11391 7262 11392
rect 790 11188 796 11252
rect 860 11250 866 11252
rect 1485 11250 1551 11253
rect 860 11248 1551 11250
rect 860 11192 1490 11248
rect 1546 11192 1551 11248
rect 860 11190 1551 11192
rect 860 11188 866 11190
rect 1485 11187 1551 11190
rect 5625 11116 5691 11117
rect 5574 11052 5580 11116
rect 5644 11114 5691 11116
rect 5644 11112 5736 11114
rect 5686 11056 5736 11112
rect 5644 11054 5736 11056
rect 5644 11052 5691 11054
rect 5625 11051 5691 11052
rect 2606 10912 2922 10913
rect 2606 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2922 10912
rect 2606 10847 2922 10848
rect 7606 10912 7922 10913
rect 7606 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7922 10912
rect 7606 10847 7922 10848
rect 3969 10842 4035 10845
rect 3969 10840 7482 10842
rect 3969 10784 3974 10840
rect 4030 10784 7482 10840
rect 3969 10782 7482 10784
rect 3969 10779 4035 10782
rect 3509 10706 3575 10709
rect 7281 10706 7347 10709
rect 3509 10704 7347 10706
rect 3509 10648 3514 10704
rect 3570 10648 7286 10704
rect 7342 10648 7347 10704
rect 3509 10646 7347 10648
rect 7422 10706 7482 10782
rect 8753 10706 8819 10709
rect 11108 10706 11908 10736
rect 7422 10646 8402 10706
rect 3509 10643 3575 10646
rect 7281 10643 7347 10646
rect 1669 10570 1735 10573
rect 8109 10570 8175 10573
rect 1669 10568 8175 10570
rect 1669 10512 1674 10568
rect 1730 10512 8114 10568
rect 8170 10512 8175 10568
rect 1669 10510 8175 10512
rect 8342 10570 8402 10646
rect 8753 10704 11908 10706
rect 8753 10648 8758 10704
rect 8814 10648 11908 10704
rect 8753 10646 11908 10648
rect 8753 10643 8819 10646
rect 11108 10616 11908 10646
rect 9121 10570 9187 10573
rect 8342 10568 9187 10570
rect 8342 10512 9126 10568
rect 9182 10512 9187 10568
rect 8342 10510 9187 10512
rect 1669 10507 1735 10510
rect 8109 10507 8175 10510
rect 9121 10507 9187 10510
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 6946 10368 7262 10369
rect 6946 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7262 10368
rect 6946 10303 7262 10304
rect 2998 10236 3004 10300
rect 3068 10298 3074 10300
rect 3141 10298 3207 10301
rect 3068 10296 3207 10298
rect 3068 10240 3146 10296
rect 3202 10240 3207 10296
rect 3068 10238 3207 10240
rect 3068 10236 3074 10238
rect 3141 10235 3207 10238
rect 3601 10298 3667 10301
rect 3601 10296 6746 10298
rect 3601 10240 3606 10296
rect 3662 10240 6746 10296
rect 3601 10238 6746 10240
rect 3601 10235 3667 10238
rect 6177 10162 6243 10165
rect 6310 10162 6316 10164
rect 6177 10160 6316 10162
rect 6177 10104 6182 10160
rect 6238 10104 6316 10160
rect 6177 10102 6316 10104
rect 6177 10099 6243 10102
rect 6310 10100 6316 10102
rect 6380 10100 6386 10164
rect 6686 10162 6746 10238
rect 9949 10162 10015 10165
rect 6686 10160 10015 10162
rect 6686 10104 9954 10160
rect 10010 10104 10015 10160
rect 6686 10102 10015 10104
rect 9949 10099 10015 10102
rect 2313 10026 2379 10029
rect 2313 10024 8218 10026
rect 2313 9968 2318 10024
rect 2374 9968 8218 10024
rect 2313 9966 8218 9968
rect 2313 9963 2379 9966
rect 4429 9890 4495 9893
rect 4654 9890 4660 9892
rect 4429 9888 4660 9890
rect 4429 9832 4434 9888
rect 4490 9832 4660 9888
rect 4429 9830 4660 9832
rect 4429 9827 4495 9830
rect 4654 9828 4660 9830
rect 4724 9828 4730 9892
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 7606 9824 7922 9825
rect 7606 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7922 9824
rect 7606 9759 7922 9760
rect 3233 9756 3299 9757
rect 3182 9692 3188 9756
rect 3252 9754 3299 9756
rect 3252 9752 3344 9754
rect 3294 9696 3344 9752
rect 3252 9694 3344 9696
rect 3252 9692 3299 9694
rect 4470 9692 4476 9756
rect 4540 9754 4546 9756
rect 5533 9754 5599 9757
rect 8158 9756 8218 9966
rect 4540 9752 5599 9754
rect 4540 9696 5538 9752
rect 5594 9696 5599 9752
rect 4540 9694 5599 9696
rect 4540 9692 4546 9694
rect 3233 9691 3299 9692
rect 5533 9691 5599 9694
rect 8150 9692 8156 9756
rect 8220 9692 8226 9756
rect 1853 9618 1919 9621
rect 10133 9618 10199 9621
rect 11108 9618 11908 9648
rect 1853 9616 8034 9618
rect 1853 9560 1858 9616
rect 1914 9560 8034 9616
rect 1853 9558 8034 9560
rect 1853 9555 1919 9558
rect 2313 9482 2379 9485
rect 7833 9482 7899 9485
rect 2313 9480 7899 9482
rect 2313 9424 2318 9480
rect 2374 9424 7838 9480
rect 7894 9424 7899 9480
rect 2313 9422 7899 9424
rect 2313 9419 2379 9422
rect 7833 9419 7899 9422
rect 7974 9346 8034 9558
rect 10133 9616 11908 9618
rect 10133 9560 10138 9616
rect 10194 9560 11908 9616
rect 10133 9558 11908 9560
rect 10133 9555 10199 9558
rect 11108 9528 11908 9558
rect 9765 9484 9831 9485
rect 9765 9482 9812 9484
rect 9720 9480 9812 9482
rect 9720 9424 9770 9480
rect 9720 9422 9812 9424
rect 9765 9420 9812 9422
rect 9876 9420 9882 9484
rect 9765 9419 9831 9420
rect 10041 9346 10107 9349
rect 7974 9344 10107 9346
rect 7974 9288 10046 9344
rect 10102 9288 10107 9344
rect 7974 9286 10107 9288
rect 10041 9283 10107 9286
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 6946 9280 7262 9281
rect 6946 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7262 9280
rect 6946 9215 7262 9216
rect 3601 9074 3667 9077
rect 8017 9074 8083 9077
rect 3601 9072 8083 9074
rect 3601 9016 3606 9072
rect 3662 9016 8022 9072
rect 8078 9016 8083 9072
rect 3601 9014 8083 9016
rect 3601 9011 3667 9014
rect 8017 9011 8083 9014
rect 2773 8938 2839 8941
rect 3550 8938 3556 8940
rect 2773 8936 3556 8938
rect 2773 8880 2778 8936
rect 2834 8880 3556 8936
rect 2773 8878 3556 8880
rect 2773 8875 2839 8878
rect 3550 8876 3556 8878
rect 3620 8876 3626 8940
rect 5206 8876 5212 8940
rect 5276 8938 5282 8940
rect 7557 8938 7623 8941
rect 5276 8936 7623 8938
rect 5276 8880 7562 8936
rect 7618 8880 7623 8936
rect 5276 8878 7623 8880
rect 5276 8876 5282 8878
rect 7557 8875 7623 8878
rect 3969 8804 4035 8805
rect 3918 8802 3924 8804
rect 3878 8742 3924 8802
rect 3988 8800 4035 8804
rect 4030 8744 4035 8800
rect 3918 8740 3924 8742
rect 3988 8740 4035 8744
rect 3969 8739 4035 8740
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 7606 8736 7922 8737
rect 7606 8672 7612 8736
rect 7676 8672 7692 8736
rect 7756 8672 7772 8736
rect 7836 8672 7852 8736
rect 7916 8672 7922 8736
rect 7606 8671 7922 8672
rect 2405 8530 2471 8533
rect 4521 8530 4587 8533
rect 2405 8528 4587 8530
rect 2405 8472 2410 8528
rect 2466 8472 4526 8528
rect 4582 8472 4587 8528
rect 2405 8470 4587 8472
rect 2405 8467 2471 8470
rect 4521 8467 4587 8470
rect 10409 8530 10475 8533
rect 11108 8530 11908 8560
rect 10409 8528 11908 8530
rect 10409 8472 10414 8528
rect 10470 8472 11908 8528
rect 10409 8470 11908 8472
rect 10409 8467 10475 8470
rect 11108 8440 11908 8470
rect 1945 8394 2011 8397
rect 5533 8394 5599 8397
rect 1945 8392 5599 8394
rect 1945 8336 1950 8392
rect 2006 8336 5538 8392
rect 5594 8336 5599 8392
rect 1945 8334 5599 8336
rect 1945 8331 2011 8334
rect 5533 8331 5599 8334
rect 3969 8258 4035 8261
rect 4102 8258 4108 8260
rect 3969 8256 4108 8258
rect 3969 8200 3974 8256
rect 4030 8200 4108 8256
rect 3969 8198 4108 8200
rect 3969 8195 4035 8198
rect 4102 8196 4108 8198
rect 4172 8196 4178 8260
rect 4337 8258 4403 8261
rect 9213 8260 9279 8261
rect 4470 8258 4476 8260
rect 4337 8256 4476 8258
rect 4337 8200 4342 8256
rect 4398 8200 4476 8256
rect 4337 8198 4476 8200
rect 4337 8195 4403 8198
rect 4470 8196 4476 8198
rect 4540 8196 4546 8260
rect 9213 8258 9260 8260
rect 9168 8256 9260 8258
rect 9168 8200 9218 8256
rect 9168 8198 9260 8200
rect 9213 8196 9260 8198
rect 9324 8196 9330 8260
rect 9213 8195 9279 8196
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 6946 8192 7262 8193
rect 6946 8128 6952 8192
rect 7016 8128 7032 8192
rect 7096 8128 7112 8192
rect 7176 8128 7192 8192
rect 7256 8128 7262 8192
rect 6946 8127 7262 8128
rect 2998 8060 3004 8124
rect 3068 8122 3074 8124
rect 5257 8122 5323 8125
rect 3068 8120 5323 8122
rect 3068 8064 5262 8120
rect 5318 8064 5323 8120
rect 3068 8062 5323 8064
rect 3068 8060 3074 8062
rect 5257 8059 5323 8062
rect 8753 8122 8819 8125
rect 9305 8122 9371 8125
rect 10409 8122 10475 8125
rect 8753 8120 10475 8122
rect 8753 8064 8758 8120
rect 8814 8064 9310 8120
rect 9366 8064 10414 8120
rect 10470 8064 10475 8120
rect 8753 8062 10475 8064
rect 8753 8059 8819 8062
rect 9305 8059 9371 8062
rect 10409 8059 10475 8062
rect 3969 7986 4035 7989
rect 6729 7986 6795 7989
rect 7414 7986 7420 7988
rect 3969 7984 7420 7986
rect 3969 7928 3974 7984
rect 4030 7928 6734 7984
rect 6790 7928 7420 7984
rect 3969 7926 7420 7928
rect 3969 7923 4035 7926
rect 6729 7923 6795 7926
rect 7414 7924 7420 7926
rect 7484 7924 7490 7988
rect 8293 7986 8359 7989
rect 10409 7986 10475 7989
rect 8293 7984 10475 7986
rect 8293 7928 8298 7984
rect 8354 7928 10414 7984
rect 10470 7928 10475 7984
rect 8293 7926 10475 7928
rect 8293 7923 8359 7926
rect 10409 7923 10475 7926
rect 6678 7788 6684 7852
rect 6748 7850 6754 7852
rect 8201 7850 8267 7853
rect 6748 7848 8267 7850
rect 6748 7792 8206 7848
rect 8262 7792 8267 7848
rect 6748 7790 8267 7792
rect 6748 7788 6754 7790
rect 8201 7787 8267 7790
rect 8753 7850 8819 7853
rect 9213 7850 9279 7853
rect 8753 7848 9279 7850
rect 8753 7792 8758 7848
rect 8814 7792 9218 7848
rect 9274 7792 9279 7848
rect 8753 7790 9279 7792
rect 8753 7787 8819 7790
rect 9213 7787 9279 7790
rect 3141 7714 3207 7717
rect 3366 7714 3372 7716
rect 3141 7712 3372 7714
rect 3141 7656 3146 7712
rect 3202 7656 3372 7712
rect 3141 7654 3372 7656
rect 3141 7651 3207 7654
rect 3366 7652 3372 7654
rect 3436 7652 3442 7716
rect 8753 7714 8819 7717
rect 9213 7714 9279 7717
rect 8753 7712 9279 7714
rect 8753 7656 8758 7712
rect 8814 7656 9218 7712
rect 9274 7656 9279 7712
rect 8753 7654 9279 7656
rect 8753 7651 8819 7654
rect 9213 7651 9279 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 7606 7583 7922 7584
rect 3693 7578 3759 7581
rect 5390 7578 5396 7580
rect 3693 7576 5396 7578
rect 3693 7520 3698 7576
rect 3754 7520 5396 7576
rect 3693 7518 5396 7520
rect 3693 7515 3759 7518
rect 5390 7516 5396 7518
rect 5460 7516 5466 7580
rect 3693 7442 3759 7445
rect 10133 7442 10199 7445
rect 3693 7440 10199 7442
rect 3693 7384 3698 7440
rect 3754 7384 10138 7440
rect 10194 7384 10199 7440
rect 3693 7382 10199 7384
rect 3693 7379 3759 7382
rect 10133 7379 10199 7382
rect 10409 7442 10475 7445
rect 11108 7442 11908 7472
rect 10409 7440 11908 7442
rect 10409 7384 10414 7440
rect 10470 7384 11908 7440
rect 10409 7382 11908 7384
rect 10409 7379 10475 7382
rect 11108 7352 11908 7382
rect 2865 7306 2931 7309
rect 6913 7306 6979 7309
rect 2865 7304 6979 7306
rect 2865 7248 2870 7304
rect 2926 7248 6918 7304
rect 6974 7248 6979 7304
rect 2865 7246 6979 7248
rect 2865 7243 2931 7246
rect 6913 7243 6979 7246
rect 2497 7170 2563 7173
rect 4705 7170 4771 7173
rect 2497 7168 4771 7170
rect 2497 7112 2502 7168
rect 2558 7112 4710 7168
rect 4766 7112 4771 7168
rect 2497 7110 4771 7112
rect 2497 7107 2563 7110
rect 4705 7107 4771 7110
rect 5758 7108 5764 7172
rect 5828 7170 5834 7172
rect 5901 7170 5967 7173
rect 10317 7170 10383 7173
rect 5828 7168 5967 7170
rect 5828 7112 5906 7168
rect 5962 7112 5967 7168
rect 5828 7110 5967 7112
rect 5828 7108 5834 7110
rect 5901 7107 5967 7110
rect 7422 7168 10383 7170
rect 7422 7112 10322 7168
rect 10378 7112 10383 7168
rect 7422 7110 10383 7112
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 3182 7034 3188 7036
rect 2730 6974 3188 7034
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 1945 6898 2011 6901
rect 2730 6898 2790 6974
rect 3182 6972 3188 6974
rect 3252 7034 3258 7036
rect 3252 6974 6746 7034
rect 3252 6972 3258 6974
rect 1945 6896 2790 6898
rect 1945 6840 1950 6896
rect 2006 6840 2790 6896
rect 1945 6838 2790 6840
rect 2865 6898 2931 6901
rect 3417 6898 3483 6901
rect 4061 6898 4127 6901
rect 5206 6898 5212 6900
rect 2865 6896 4127 6898
rect 2865 6840 2870 6896
rect 2926 6840 3422 6896
rect 3478 6840 4066 6896
rect 4122 6840 4127 6896
rect 2865 6838 4127 6840
rect 1945 6835 2011 6838
rect 2865 6835 2931 6838
rect 3417 6835 3483 6838
rect 4061 6835 4127 6838
rect 4432 6838 5212 6898
rect 2681 6762 2747 6765
rect 4432 6762 4492 6838
rect 5206 6836 5212 6838
rect 5276 6836 5282 6900
rect 6269 6898 6335 6901
rect 6494 6898 6500 6900
rect 6269 6896 6500 6898
rect 6269 6840 6274 6896
rect 6330 6840 6500 6896
rect 6269 6838 6500 6840
rect 6269 6835 6335 6838
rect 6494 6836 6500 6838
rect 6564 6836 6570 6900
rect 6686 6898 6746 6974
rect 7422 6898 7482 7110
rect 10317 7107 10383 7110
rect 6686 6838 7482 6898
rect 7557 6898 7623 6901
rect 9806 6898 9812 6900
rect 7557 6896 9812 6898
rect 7557 6840 7562 6896
rect 7618 6840 9812 6896
rect 7557 6838 9812 6840
rect 7557 6835 7623 6838
rect 9806 6836 9812 6838
rect 9876 6898 9882 6900
rect 10317 6898 10383 6901
rect 9876 6896 10383 6898
rect 9876 6840 10322 6896
rect 10378 6840 10383 6896
rect 9876 6838 10383 6840
rect 9876 6836 9882 6838
rect 10317 6835 10383 6838
rect 2681 6760 4492 6762
rect 2681 6704 2686 6760
rect 2742 6704 4492 6760
rect 2681 6702 4492 6704
rect 2681 6699 2747 6702
rect 6310 6700 6316 6764
rect 6380 6762 6386 6764
rect 6380 6702 8586 6762
rect 6380 6700 6386 6702
rect 4889 6626 4955 6629
rect 6821 6626 6887 6629
rect 8526 6628 8586 6702
rect 4889 6624 6887 6626
rect 4889 6568 4894 6624
rect 4950 6568 6826 6624
rect 6882 6568 6887 6624
rect 4889 6566 6887 6568
rect 4889 6563 4955 6566
rect 6821 6563 6887 6566
rect 8518 6564 8524 6628
rect 8588 6626 8594 6628
rect 8661 6626 8727 6629
rect 8588 6624 8727 6626
rect 8588 6568 8666 6624
rect 8722 6568 8727 6624
rect 8588 6566 8727 6568
rect 8588 6564 8594 6566
rect 8661 6563 8727 6566
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 7606 6495 7922 6496
rect 5717 6490 5783 6493
rect 6913 6490 6979 6493
rect 5717 6488 6979 6490
rect 5717 6432 5722 6488
rect 5778 6432 6918 6488
rect 6974 6432 6979 6488
rect 5717 6430 6979 6432
rect 5717 6427 5783 6430
rect 6913 6427 6979 6430
rect 2681 6354 2747 6357
rect 2998 6354 3004 6356
rect 2681 6352 3004 6354
rect 2681 6296 2686 6352
rect 2742 6296 3004 6352
rect 2681 6294 3004 6296
rect 2681 6291 2747 6294
rect 2998 6292 3004 6294
rect 3068 6292 3074 6356
rect 4654 6292 4660 6356
rect 4724 6354 4730 6356
rect 4889 6354 4955 6357
rect 8661 6354 8727 6357
rect 4724 6352 8727 6354
rect 4724 6296 4894 6352
rect 4950 6296 8666 6352
rect 8722 6296 8727 6352
rect 4724 6294 8727 6296
rect 4724 6292 4730 6294
rect 4889 6291 4955 6294
rect 8661 6291 8727 6294
rect 10409 6354 10475 6357
rect 11108 6354 11908 6384
rect 10409 6352 11908 6354
rect 10409 6296 10414 6352
rect 10470 6296 11908 6352
rect 10409 6294 11908 6296
rect 10409 6291 10475 6294
rect 11108 6264 11908 6294
rect 2221 6218 2287 6221
rect 6637 6218 6703 6221
rect 2221 6216 6703 6218
rect 2221 6160 2226 6216
rect 2282 6160 6642 6216
rect 6698 6160 6703 6216
rect 2221 6158 6703 6160
rect 2221 6155 2287 6158
rect 6637 6155 6703 6158
rect 6821 6218 6887 6221
rect 9213 6220 9279 6221
rect 9213 6218 9260 6220
rect 6821 6216 9260 6218
rect 6821 6160 6826 6216
rect 6882 6160 9218 6216
rect 6821 6158 9260 6160
rect 6821 6155 6887 6158
rect 9213 6156 9260 6158
rect 9324 6156 9330 6220
rect 9397 6216 9463 6221
rect 9397 6160 9402 6216
rect 9458 6160 9463 6216
rect 9213 6155 9279 6156
rect 9397 6155 9463 6160
rect 3509 6082 3575 6085
rect 6637 6082 6703 6085
rect 3509 6080 6703 6082
rect 3509 6024 3514 6080
rect 3570 6024 6642 6080
rect 6698 6024 6703 6080
rect 3509 6022 6703 6024
rect 3509 6019 3575 6022
rect 6637 6019 6703 6022
rect 8477 6082 8543 6085
rect 9400 6082 9460 6155
rect 8477 6080 9460 6082
rect 8477 6024 8482 6080
rect 8538 6024 9460 6080
rect 8477 6022 9460 6024
rect 8477 6019 8543 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 3141 5946 3207 5949
rect 2454 5944 3207 5946
rect 2454 5888 3146 5944
rect 3202 5888 3207 5944
rect 2454 5886 3207 5888
rect 2221 5810 2287 5813
rect 2454 5810 2514 5886
rect 3141 5883 3207 5886
rect 3969 5946 4035 5949
rect 6269 5946 6335 5949
rect 3969 5944 6335 5946
rect 3969 5888 3974 5944
rect 4030 5888 6274 5944
rect 6330 5888 6335 5944
rect 3969 5886 6335 5888
rect 3969 5883 4035 5886
rect 6269 5883 6335 5886
rect 2221 5808 2514 5810
rect 2221 5752 2226 5808
rect 2282 5752 2514 5808
rect 2221 5750 2514 5752
rect 2589 5810 2655 5813
rect 10225 5810 10291 5813
rect 2589 5808 10291 5810
rect 2589 5752 2594 5808
rect 2650 5752 10230 5808
rect 10286 5752 10291 5808
rect 2589 5750 10291 5752
rect 2221 5747 2287 5750
rect 2589 5747 2655 5750
rect 10225 5747 10291 5750
rect 1025 5674 1091 5677
rect 5441 5674 5507 5677
rect 1025 5672 5507 5674
rect 1025 5616 1030 5672
rect 1086 5616 5446 5672
rect 5502 5616 5507 5672
rect 1025 5614 5507 5616
rect 1025 5611 1091 5614
rect 5441 5611 5507 5614
rect 5717 5674 5783 5677
rect 8477 5674 8543 5677
rect 5717 5672 8543 5674
rect 5717 5616 5722 5672
rect 5778 5616 8482 5672
rect 8538 5616 8543 5672
rect 5717 5614 8543 5616
rect 5717 5611 5783 5614
rect 8477 5611 8543 5614
rect 8661 5674 8727 5677
rect 9213 5674 9279 5677
rect 8661 5672 9279 5674
rect 8661 5616 8666 5672
rect 8722 5616 9218 5672
rect 9274 5616 9279 5672
rect 8661 5614 9279 5616
rect 8661 5611 8727 5614
rect 9213 5611 9279 5614
rect 3325 5538 3391 5541
rect 5625 5538 5691 5541
rect 3325 5536 5691 5538
rect 3325 5480 3330 5536
rect 3386 5480 5630 5536
rect 5686 5480 5691 5536
rect 3325 5478 5691 5480
rect 3325 5475 3391 5478
rect 5625 5475 5691 5478
rect 6269 5538 6335 5541
rect 6729 5540 6795 5541
rect 8201 5540 8267 5541
rect 6494 5538 6500 5540
rect 6269 5536 6500 5538
rect 6269 5480 6274 5536
rect 6330 5480 6500 5536
rect 6269 5478 6500 5480
rect 6269 5475 6335 5478
rect 6494 5476 6500 5478
rect 6564 5476 6570 5540
rect 6678 5476 6684 5540
rect 6748 5538 6795 5540
rect 8150 5538 8156 5540
rect 6748 5536 6840 5538
rect 6790 5480 6840 5536
rect 6748 5478 6840 5480
rect 8110 5478 8156 5538
rect 8220 5536 8267 5540
rect 8262 5480 8267 5536
rect 6748 5476 6795 5478
rect 8150 5476 8156 5478
rect 8220 5476 8267 5480
rect 6729 5475 6795 5476
rect 8201 5475 8267 5476
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 7606 5407 7922 5408
rect 3325 5402 3391 5405
rect 3918 5402 3924 5404
rect 3325 5400 3924 5402
rect 3325 5344 3330 5400
rect 3386 5344 3924 5400
rect 3325 5342 3924 5344
rect 3325 5339 3391 5342
rect 3918 5340 3924 5342
rect 3988 5340 3994 5404
rect 4102 5340 4108 5404
rect 4172 5402 4178 5404
rect 4705 5402 4771 5405
rect 4172 5400 4771 5402
rect 4172 5344 4710 5400
rect 4766 5344 4771 5400
rect 4172 5342 4771 5344
rect 4172 5340 4178 5342
rect 4705 5339 4771 5342
rect 5574 5340 5580 5404
rect 5644 5402 5650 5404
rect 5809 5402 5875 5405
rect 5644 5400 5875 5402
rect 5644 5344 5814 5400
rect 5870 5344 5875 5400
rect 5644 5342 5875 5344
rect 5644 5340 5650 5342
rect 5809 5339 5875 5342
rect 1945 5266 2011 5269
rect 8293 5266 8359 5269
rect 1945 5264 8359 5266
rect 1945 5208 1950 5264
rect 2006 5208 8298 5264
rect 8354 5208 8359 5264
rect 1945 5206 8359 5208
rect 1945 5203 2011 5206
rect 8293 5203 8359 5206
rect 10409 5266 10475 5269
rect 11108 5266 11908 5296
rect 10409 5264 11908 5266
rect 10409 5208 10414 5264
rect 10470 5208 11908 5264
rect 10409 5206 11908 5208
rect 10409 5203 10475 5206
rect 11108 5176 11908 5206
rect 3049 5130 3115 5133
rect 8201 5130 8267 5133
rect 3049 5128 8267 5130
rect 3049 5072 3054 5128
rect 3110 5072 8206 5128
rect 8262 5072 8267 5128
rect 3049 5070 8267 5072
rect 3049 5067 3115 5070
rect 8201 5067 8267 5070
rect 3141 4994 3207 4997
rect 3366 4994 3372 4996
rect 3141 4992 3372 4994
rect 3141 4936 3146 4992
rect 3202 4936 3372 4992
rect 3141 4934 3372 4936
rect 3141 4931 3207 4934
rect 3366 4932 3372 4934
rect 3436 4994 3442 4996
rect 6729 4994 6795 4997
rect 3436 4992 6795 4994
rect 3436 4936 6734 4992
rect 6790 4936 6795 4992
rect 3436 4934 6795 4936
rect 3436 4932 3442 4934
rect 6729 4931 6795 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 3877 4858 3943 4861
rect 6545 4858 6611 4861
rect 3877 4856 6611 4858
rect 3877 4800 3882 4856
rect 3938 4800 6550 4856
rect 6606 4800 6611 4856
rect 3877 4798 6611 4800
rect 3877 4795 3943 4798
rect 6545 4795 6611 4798
rect 1301 4722 1367 4725
rect 9949 4722 10015 4725
rect 1301 4720 10015 4722
rect 1301 4664 1306 4720
rect 1362 4664 9954 4720
rect 10010 4664 10015 4720
rect 1301 4662 10015 4664
rect 1301 4659 1367 4662
rect 9949 4659 10015 4662
rect 5165 4586 5231 4589
rect 9581 4586 9647 4589
rect 5165 4584 9647 4586
rect 5165 4528 5170 4584
rect 5226 4528 9586 4584
rect 9642 4528 9647 4584
rect 5165 4526 9647 4528
rect 5165 4523 5231 4526
rect 9581 4523 9647 4526
rect 4889 4450 4955 4453
rect 6821 4450 6887 4453
rect 4889 4448 6887 4450
rect 4889 4392 4894 4448
rect 4950 4392 6826 4448
rect 6882 4392 6887 4448
rect 4889 4390 6887 4392
rect 4889 4387 4955 4390
rect 6821 4387 6887 4390
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 7606 4319 7922 4320
rect 5349 4316 5415 4317
rect 5349 4312 5396 4316
rect 5460 4314 5466 4316
rect 5349 4256 5354 4312
rect 5349 4252 5396 4256
rect 5460 4254 5506 4314
rect 5460 4252 5466 4254
rect 5349 4251 5415 4252
rect 1853 4178 1919 4181
rect 5901 4178 5967 4181
rect 1853 4176 5967 4178
rect 1853 4120 1858 4176
rect 1914 4120 5906 4176
rect 5962 4120 5967 4176
rect 1853 4118 5967 4120
rect 1853 4115 1919 4118
rect 5901 4115 5967 4118
rect 7414 4116 7420 4180
rect 7484 4178 7490 4180
rect 7833 4178 7899 4181
rect 7484 4176 7899 4178
rect 7484 4120 7838 4176
rect 7894 4120 7899 4176
rect 7484 4118 7899 4120
rect 7484 4116 7490 4118
rect 7833 4115 7899 4118
rect 10409 4178 10475 4181
rect 11108 4178 11908 4208
rect 10409 4176 11908 4178
rect 10409 4120 10414 4176
rect 10470 4120 11908 4176
rect 10409 4118 11908 4120
rect 10409 4115 10475 4118
rect 11108 4088 11908 4118
rect 1117 4042 1183 4045
rect 9397 4042 9463 4045
rect 1117 4040 9463 4042
rect 1117 3984 1122 4040
rect 1178 3984 9402 4040
rect 9458 3984 9463 4040
rect 1117 3982 9463 3984
rect 1117 3979 1183 3982
rect 9397 3979 9463 3982
rect 5809 3908 5875 3909
rect 5758 3844 5764 3908
rect 5828 3906 5875 3908
rect 5828 3904 5920 3906
rect 5870 3848 5920 3904
rect 5828 3846 5920 3848
rect 5828 3844 5875 3846
rect 5809 3843 5875 3844
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 5206 3708 5212 3772
rect 5276 3770 5282 3772
rect 5533 3770 5599 3773
rect 5276 3768 5599 3770
rect 5276 3712 5538 3768
rect 5594 3712 5599 3768
rect 5276 3710 5599 3712
rect 5276 3708 5282 3710
rect 5533 3707 5599 3710
rect 2037 3634 2103 3637
rect 9213 3634 9279 3637
rect 2037 3632 9279 3634
rect 2037 3576 2042 3632
rect 2098 3576 9218 3632
rect 9274 3576 9279 3632
rect 2037 3574 9279 3576
rect 2037 3571 2103 3574
rect 9213 3571 9279 3574
rect 4153 3498 4219 3501
rect 8518 3498 8524 3500
rect 4153 3496 8524 3498
rect 4153 3440 4158 3496
rect 4214 3440 8524 3496
rect 4153 3438 8524 3440
rect 4153 3435 4219 3438
rect 8518 3436 8524 3438
rect 8588 3436 8594 3500
rect 3550 3300 3556 3364
rect 3620 3362 3626 3364
rect 4705 3362 4771 3365
rect 3620 3360 4771 3362
rect 3620 3304 4710 3360
rect 4766 3304 4771 3360
rect 3620 3302 4771 3304
rect 3620 3300 3626 3302
rect 4705 3299 4771 3302
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 7606 3231 7922 3232
rect 10409 3090 10475 3093
rect 11108 3090 11908 3120
rect 10409 3088 11908 3090
rect 10409 3032 10414 3088
rect 10470 3032 11908 3088
rect 10409 3030 11908 3032
rect 10409 3027 10475 3030
rect 11108 3000 11908 3030
rect 2957 2954 3023 2957
rect 4061 2954 4127 2957
rect 10317 2954 10383 2957
rect 2957 2952 10383 2954
rect 2957 2896 2962 2952
rect 3018 2896 4066 2952
rect 4122 2896 10322 2952
rect 10378 2896 10383 2952
rect 2957 2894 10383 2896
rect 2957 2891 3023 2894
rect 4061 2891 4127 2894
rect 10317 2891 10383 2894
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 6946 2687 7262 2688
rect 0 2274 800 2304
rect 1025 2274 1091 2277
rect 0 2272 1091 2274
rect 0 2216 1030 2272
rect 1086 2216 1091 2272
rect 0 2214 1091 2216
rect 0 2184 800 2214
rect 1025 2211 1091 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 7606 2143 7922 2144
rect 10133 2002 10199 2005
rect 11108 2002 11908 2032
rect 10133 2000 11908 2002
rect 10133 1944 10138 2000
rect 10194 1944 11908 2000
rect 10133 1942 11908 1944
rect 10133 1939 10199 1942
rect 11108 1912 11908 1942
rect 10869 914 10935 917
rect 11108 914 11908 944
rect 10869 912 11908 914
rect 10869 856 10874 912
rect 10930 856 11908 912
rect 10869 854 11908 856
rect 10869 851 10935 854
rect 11108 824 11908 854
<< via3 >>
rect 796 11460 860 11524
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 6952 11452 7016 11456
rect 6952 11396 6956 11452
rect 6956 11396 7012 11452
rect 7012 11396 7016 11452
rect 6952 11392 7016 11396
rect 7032 11452 7096 11456
rect 7032 11396 7036 11452
rect 7036 11396 7092 11452
rect 7092 11396 7096 11452
rect 7032 11392 7096 11396
rect 7112 11452 7176 11456
rect 7112 11396 7116 11452
rect 7116 11396 7172 11452
rect 7172 11396 7176 11452
rect 7112 11392 7176 11396
rect 7192 11452 7256 11456
rect 7192 11396 7196 11452
rect 7196 11396 7252 11452
rect 7252 11396 7256 11452
rect 7192 11392 7256 11396
rect 796 11188 860 11252
rect 5580 11112 5644 11116
rect 5580 11056 5630 11112
rect 5630 11056 5644 11112
rect 5580 11052 5644 11056
rect 2612 10908 2676 10912
rect 2612 10852 2616 10908
rect 2616 10852 2672 10908
rect 2672 10852 2676 10908
rect 2612 10848 2676 10852
rect 2692 10908 2756 10912
rect 2692 10852 2696 10908
rect 2696 10852 2752 10908
rect 2752 10852 2756 10908
rect 2692 10848 2756 10852
rect 2772 10908 2836 10912
rect 2772 10852 2776 10908
rect 2776 10852 2832 10908
rect 2832 10852 2836 10908
rect 2772 10848 2836 10852
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 7612 10908 7676 10912
rect 7612 10852 7616 10908
rect 7616 10852 7672 10908
rect 7672 10852 7676 10908
rect 7612 10848 7676 10852
rect 7692 10908 7756 10912
rect 7692 10852 7696 10908
rect 7696 10852 7752 10908
rect 7752 10852 7756 10908
rect 7692 10848 7756 10852
rect 7772 10908 7836 10912
rect 7772 10852 7776 10908
rect 7776 10852 7832 10908
rect 7832 10852 7836 10908
rect 7772 10848 7836 10852
rect 7852 10908 7916 10912
rect 7852 10852 7856 10908
rect 7856 10852 7912 10908
rect 7912 10852 7916 10908
rect 7852 10848 7916 10852
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 6952 10364 7016 10368
rect 6952 10308 6956 10364
rect 6956 10308 7012 10364
rect 7012 10308 7016 10364
rect 6952 10304 7016 10308
rect 7032 10364 7096 10368
rect 7032 10308 7036 10364
rect 7036 10308 7092 10364
rect 7092 10308 7096 10364
rect 7032 10304 7096 10308
rect 7112 10364 7176 10368
rect 7112 10308 7116 10364
rect 7116 10308 7172 10364
rect 7172 10308 7176 10364
rect 7112 10304 7176 10308
rect 7192 10364 7256 10368
rect 7192 10308 7196 10364
rect 7196 10308 7252 10364
rect 7252 10308 7256 10364
rect 7192 10304 7256 10308
rect 3004 10236 3068 10300
rect 6316 10100 6380 10164
rect 4660 9828 4724 9892
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 7612 9820 7676 9824
rect 7612 9764 7616 9820
rect 7616 9764 7672 9820
rect 7672 9764 7676 9820
rect 7612 9760 7676 9764
rect 7692 9820 7756 9824
rect 7692 9764 7696 9820
rect 7696 9764 7752 9820
rect 7752 9764 7756 9820
rect 7692 9760 7756 9764
rect 7772 9820 7836 9824
rect 7772 9764 7776 9820
rect 7776 9764 7832 9820
rect 7832 9764 7836 9820
rect 7772 9760 7836 9764
rect 7852 9820 7916 9824
rect 7852 9764 7856 9820
rect 7856 9764 7912 9820
rect 7912 9764 7916 9820
rect 7852 9760 7916 9764
rect 3188 9752 3252 9756
rect 3188 9696 3238 9752
rect 3238 9696 3252 9752
rect 3188 9692 3252 9696
rect 4476 9692 4540 9756
rect 8156 9692 8220 9756
rect 9812 9480 9876 9484
rect 9812 9424 9826 9480
rect 9826 9424 9876 9480
rect 9812 9420 9876 9424
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 6952 9276 7016 9280
rect 6952 9220 6956 9276
rect 6956 9220 7012 9276
rect 7012 9220 7016 9276
rect 6952 9216 7016 9220
rect 7032 9276 7096 9280
rect 7032 9220 7036 9276
rect 7036 9220 7092 9276
rect 7092 9220 7096 9276
rect 7032 9216 7096 9220
rect 7112 9276 7176 9280
rect 7112 9220 7116 9276
rect 7116 9220 7172 9276
rect 7172 9220 7176 9276
rect 7112 9216 7176 9220
rect 7192 9276 7256 9280
rect 7192 9220 7196 9276
rect 7196 9220 7252 9276
rect 7252 9220 7256 9276
rect 7192 9216 7256 9220
rect 3556 8876 3620 8940
rect 5212 8876 5276 8940
rect 3924 8800 3988 8804
rect 3924 8744 3974 8800
rect 3974 8744 3988 8800
rect 3924 8740 3988 8744
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 7612 8732 7676 8736
rect 7612 8676 7616 8732
rect 7616 8676 7672 8732
rect 7672 8676 7676 8732
rect 7612 8672 7676 8676
rect 7692 8732 7756 8736
rect 7692 8676 7696 8732
rect 7696 8676 7752 8732
rect 7752 8676 7756 8732
rect 7692 8672 7756 8676
rect 7772 8732 7836 8736
rect 7772 8676 7776 8732
rect 7776 8676 7832 8732
rect 7832 8676 7836 8732
rect 7772 8672 7836 8676
rect 7852 8732 7916 8736
rect 7852 8676 7856 8732
rect 7856 8676 7912 8732
rect 7912 8676 7916 8732
rect 7852 8672 7916 8676
rect 4108 8196 4172 8260
rect 4476 8196 4540 8260
rect 9260 8256 9324 8260
rect 9260 8200 9274 8256
rect 9274 8200 9324 8256
rect 9260 8196 9324 8200
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 6952 8188 7016 8192
rect 6952 8132 6956 8188
rect 6956 8132 7012 8188
rect 7012 8132 7016 8188
rect 6952 8128 7016 8132
rect 7032 8188 7096 8192
rect 7032 8132 7036 8188
rect 7036 8132 7092 8188
rect 7092 8132 7096 8188
rect 7032 8128 7096 8132
rect 7112 8188 7176 8192
rect 7112 8132 7116 8188
rect 7116 8132 7172 8188
rect 7172 8132 7176 8188
rect 7112 8128 7176 8132
rect 7192 8188 7256 8192
rect 7192 8132 7196 8188
rect 7196 8132 7252 8188
rect 7252 8132 7256 8188
rect 7192 8128 7256 8132
rect 3004 8060 3068 8124
rect 7420 7924 7484 7988
rect 6684 7788 6748 7852
rect 3372 7652 3436 7716
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 5396 7516 5460 7580
rect 5764 7108 5828 7172
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 3188 6972 3252 7036
rect 5212 6836 5276 6900
rect 6500 6836 6564 6900
rect 9812 6836 9876 6900
rect 6316 6700 6380 6764
rect 8524 6564 8588 6628
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 3004 6292 3068 6356
rect 4660 6292 4724 6356
rect 9260 6216 9324 6220
rect 9260 6160 9274 6216
rect 9274 6160 9324 6216
rect 9260 6156 9324 6160
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 6500 5476 6564 5540
rect 6684 5536 6748 5540
rect 6684 5480 6734 5536
rect 6734 5480 6748 5536
rect 6684 5476 6748 5480
rect 8156 5536 8220 5540
rect 8156 5480 8206 5536
rect 8206 5480 8220 5536
rect 8156 5476 8220 5480
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 3924 5340 3988 5404
rect 4108 5340 4172 5404
rect 5580 5340 5644 5404
rect 3372 4932 3436 4996
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 5396 4312 5460 4316
rect 5396 4256 5410 4312
rect 5410 4256 5460 4312
rect 5396 4252 5460 4256
rect 7420 4116 7484 4180
rect 5764 3904 5828 3908
rect 5764 3848 5814 3904
rect 5814 3848 5828 3904
rect 5764 3844 5828 3848
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 5212 3708 5276 3772
rect 8524 3436 8588 3500
rect 3556 3300 3620 3364
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
<< metal4 >>
rect 795 11524 861 11525
rect 795 11460 796 11524
rect 860 11460 861 11524
rect 795 11459 861 11460
rect 798 11253 858 11459
rect 1944 11456 2264 11472
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 795 11252 861 11253
rect 795 11188 796 11252
rect 860 11188 861 11252
rect 795 11187 861 11188
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8294 2264 9216
rect 1944 8192 1986 8294
rect 2222 8192 2264 8294
rect 1944 8128 1952 8192
rect 2256 8128 2264 8192
rect 1944 8058 1986 8128
rect 2222 8058 2264 8128
rect 1944 7104 2264 8058
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 10912 2924 11472
rect 6944 11456 7264 11472
rect 6944 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7264 11456
rect 5579 11116 5645 11117
rect 5579 11052 5580 11116
rect 5644 11052 5645 11116
rect 5579 11051 5645 11052
rect 2604 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2924 10912
rect 2604 9824 2924 10848
rect 3003 10300 3069 10301
rect 3003 10236 3004 10300
rect 3068 10236 3069 10300
rect 3003 10235 3069 10236
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8954 2924 9760
rect 2604 8736 2646 8954
rect 2882 8736 2924 8954
rect 2604 8672 2612 8736
rect 2676 8672 2692 8718
rect 2756 8672 2772 8718
rect 2836 8672 2852 8718
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 3006 8125 3066 10235
rect 4659 9892 4725 9893
rect 4659 9828 4660 9892
rect 4724 9828 4725 9892
rect 4659 9827 4725 9828
rect 3187 9756 3253 9757
rect 3187 9692 3188 9756
rect 3252 9692 3253 9756
rect 3187 9691 3253 9692
rect 4475 9756 4541 9757
rect 4475 9692 4476 9756
rect 4540 9692 4541 9756
rect 4475 9691 4541 9692
rect 3003 8124 3069 8125
rect 3003 8060 3004 8124
rect 3068 8060 3069 8124
rect 3003 8059 3069 8060
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 3006 6357 3066 8059
rect 3190 7037 3250 9691
rect 3555 8940 3621 8941
rect 3555 8876 3556 8940
rect 3620 8876 3621 8940
rect 3555 8875 3621 8876
rect 3371 7716 3437 7717
rect 3371 7652 3372 7716
rect 3436 7652 3437 7716
rect 3371 7651 3437 7652
rect 3187 7036 3253 7037
rect 3187 6972 3188 7036
rect 3252 6972 3253 7036
rect 3187 6971 3253 6972
rect 3003 6356 3069 6357
rect 3003 6292 3004 6356
rect 3068 6292 3069 6356
rect 3003 6291 3069 6292
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 3374 4997 3434 7651
rect 3371 4996 3437 4997
rect 3371 4932 3372 4996
rect 3436 4932 3437 4996
rect 3371 4931 3437 4932
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 3558 3365 3618 8875
rect 3923 8804 3989 8805
rect 3923 8740 3924 8804
rect 3988 8740 3989 8804
rect 3923 8739 3989 8740
rect 3926 5405 3986 8739
rect 4478 8261 4538 9691
rect 4107 8260 4173 8261
rect 4107 8196 4108 8260
rect 4172 8196 4173 8260
rect 4107 8195 4173 8196
rect 4475 8260 4541 8261
rect 4475 8196 4476 8260
rect 4540 8196 4541 8260
rect 4475 8195 4541 8196
rect 4110 5405 4170 8195
rect 4662 6357 4722 9827
rect 5211 8940 5277 8941
rect 5211 8876 5212 8940
rect 5276 8876 5277 8940
rect 5211 8875 5277 8876
rect 5214 6901 5274 8875
rect 5395 7580 5461 7581
rect 5395 7516 5396 7580
rect 5460 7516 5461 7580
rect 5395 7515 5461 7516
rect 5211 6900 5277 6901
rect 5211 6836 5212 6900
rect 5276 6836 5277 6900
rect 5211 6835 5277 6836
rect 4659 6356 4725 6357
rect 4659 6292 4660 6356
rect 4724 6292 4725 6356
rect 4659 6291 4725 6292
rect 3923 5404 3989 5405
rect 3923 5340 3924 5404
rect 3988 5340 3989 5404
rect 3923 5339 3989 5340
rect 4107 5404 4173 5405
rect 4107 5340 4108 5404
rect 4172 5340 4173 5404
rect 4107 5339 4173 5340
rect 5214 3773 5274 6835
rect 5398 4317 5458 7515
rect 5582 5405 5642 11051
rect 6944 10368 7264 11392
rect 6944 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7264 10368
rect 6315 10164 6381 10165
rect 6315 10100 6316 10164
rect 6380 10100 6381 10164
rect 6315 10099 6381 10100
rect 5763 7172 5829 7173
rect 5763 7108 5764 7172
rect 5828 7108 5829 7172
rect 5763 7107 5829 7108
rect 5579 5404 5645 5405
rect 5579 5340 5580 5404
rect 5644 5340 5645 5404
rect 5579 5339 5645 5340
rect 5395 4316 5461 4317
rect 5395 4252 5396 4316
rect 5460 4252 5461 4316
rect 5395 4251 5461 4252
rect 5766 3909 5826 7107
rect 6318 6765 6378 10099
rect 6944 9280 7264 10304
rect 6944 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7264 9280
rect 6944 8294 7264 9216
rect 6944 8192 6986 8294
rect 7222 8192 7264 8294
rect 6944 8128 6952 8192
rect 7256 8128 7264 8192
rect 6944 8058 6986 8128
rect 7222 8058 7264 8128
rect 6683 7852 6749 7853
rect 6683 7788 6684 7852
rect 6748 7788 6749 7852
rect 6683 7787 6749 7788
rect 6499 6900 6565 6901
rect 6499 6836 6500 6900
rect 6564 6836 6565 6900
rect 6499 6835 6565 6836
rect 6315 6764 6381 6765
rect 6315 6700 6316 6764
rect 6380 6700 6381 6764
rect 6315 6699 6381 6700
rect 6502 5541 6562 6835
rect 6686 5541 6746 7787
rect 6944 7104 7264 8058
rect 7604 10912 7924 11472
rect 7604 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7924 10912
rect 7604 9824 7924 10848
rect 7604 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7924 9824
rect 7604 8954 7924 9760
rect 8155 9756 8221 9757
rect 8155 9692 8156 9756
rect 8220 9692 8221 9756
rect 8155 9691 8221 9692
rect 7604 8736 7646 8954
rect 7882 8736 7924 8954
rect 7604 8672 7612 8736
rect 7676 8672 7692 8718
rect 7756 8672 7772 8718
rect 7836 8672 7852 8718
rect 7916 8672 7924 8736
rect 7419 7988 7485 7989
rect 7419 7924 7420 7988
rect 7484 7924 7485 7988
rect 7419 7923 7485 7924
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6944 6016 7264 7040
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6499 5540 6565 5541
rect 6499 5476 6500 5540
rect 6564 5476 6565 5540
rect 6499 5475 6565 5476
rect 6683 5540 6749 5541
rect 6683 5476 6684 5540
rect 6748 5476 6749 5540
rect 6683 5475 6749 5476
rect 6944 4928 7264 5952
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 5763 3908 5829 3909
rect 5763 3844 5764 3908
rect 5828 3844 5829 3908
rect 5763 3843 5829 3844
rect 6944 3840 7264 4864
rect 7422 4181 7482 7923
rect 7604 7648 7924 8672
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7604 6560 7924 7584
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7604 5472 7924 6496
rect 8158 5541 8218 9691
rect 9811 9484 9877 9485
rect 9811 9420 9812 9484
rect 9876 9420 9877 9484
rect 9811 9419 9877 9420
rect 9259 8260 9325 8261
rect 9259 8196 9260 8260
rect 9324 8196 9325 8260
rect 9259 8195 9325 8196
rect 8523 6628 8589 6629
rect 8523 6564 8524 6628
rect 8588 6564 8589 6628
rect 8523 6563 8589 6564
rect 8155 5540 8221 5541
rect 8155 5476 8156 5540
rect 8220 5476 8221 5540
rect 8155 5475 8221 5476
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7604 4384 7924 5408
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7419 4180 7485 4181
rect 7419 4116 7420 4180
rect 7484 4116 7485 4180
rect 7419 4115 7485 4116
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 5211 3772 5277 3773
rect 5211 3708 5212 3772
rect 5276 3708 5277 3772
rect 5211 3707 5277 3708
rect 3555 3364 3621 3365
rect 3555 3300 3556 3364
rect 3620 3300 3621 3364
rect 3555 3299 3621 3300
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 6944 2128 7264 2688
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 8526 3501 8586 6563
rect 9262 6221 9322 8195
rect 9814 6901 9874 9419
rect 9811 6900 9877 6901
rect 9811 6836 9812 6900
rect 9876 6836 9877 6900
rect 9811 6835 9877 6836
rect 9259 6220 9325 6221
rect 9259 6156 9260 6220
rect 9324 6156 9325 6220
rect 9259 6155 9325 6156
rect 8523 3500 8589 3501
rect 8523 3436 8524 3500
rect 8588 3436 8589 3500
rect 8523 3435 8589 3436
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
<< via4 >>
rect 1986 8192 2222 8294
rect 1986 8128 2016 8192
rect 2016 8128 2032 8192
rect 2032 8128 2096 8192
rect 2096 8128 2112 8192
rect 2112 8128 2176 8192
rect 2176 8128 2192 8192
rect 2192 8128 2222 8192
rect 1986 8058 2222 8128
rect 1986 3058 2222 3294
rect 2646 8736 2882 8954
rect 2646 8718 2676 8736
rect 2676 8718 2692 8736
rect 2692 8718 2756 8736
rect 2756 8718 2772 8736
rect 2772 8718 2836 8736
rect 2836 8718 2852 8736
rect 2852 8718 2882 8736
rect 2646 3718 2882 3954
rect 6986 8192 7222 8294
rect 6986 8128 7016 8192
rect 7016 8128 7032 8192
rect 7032 8128 7096 8192
rect 7096 8128 7112 8192
rect 7112 8128 7176 8192
rect 7176 8128 7192 8192
rect 7192 8128 7222 8192
rect 6986 8058 7222 8128
rect 7646 8736 7882 8954
rect 7646 8718 7676 8736
rect 7676 8718 7692 8736
rect 7692 8718 7756 8736
rect 7756 8718 7772 8736
rect 7772 8718 7836 8736
rect 7836 8718 7852 8736
rect 7852 8718 7882 8736
rect 6986 3058 7222 3294
rect 7646 3718 7882 3954
<< metal5 >>
rect 1056 8954 10812 8996
rect 1056 8718 2646 8954
rect 2882 8718 7646 8954
rect 7882 8718 10812 8954
rect 1056 8676 10812 8718
rect 1056 8294 10812 8336
rect 1056 8058 1986 8294
rect 2222 8058 6986 8294
rect 7222 8058 10812 8294
rect 1056 8016 10812 8058
rect 1056 3954 10812 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 10812 3954
rect 1056 3676 10812 3718
rect 1056 3294 10812 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 10812 3294
rect 1056 3016 10812 3058
use sky130_fd_sc_hd__and4_1  _094_
timestamp 1713593032
transform 1 0 8556 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _095_
timestamp 1713593032
transform 1 0 1472 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _096_
timestamp 1713593032
transform 1 0 3220 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _097_
timestamp 1713593032
transform -1 0 10304 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _098_
timestamp 1713593032
transform -1 0 6164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1713593032
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _100_
timestamp 1713593032
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1713593032
transform -1 0 8464 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _102_
timestamp 1713593032
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _103_
timestamp 1713593032
transform 1 0 8556 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _104_
timestamp 1713593032
transform -1 0 10304 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1713593032
transform 1 0 9476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _106_
timestamp 1713593032
transform -1 0 6256 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _107_
timestamp 1713593032
transform -1 0 9660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _108_
timestamp 1713593032
transform 1 0 2668 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1713593032
transform -1 0 6348 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _110_
timestamp 1713593032
transform -1 0 4692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _111_
timestamp 1713593032
transform 1 0 2392 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _112_
timestamp 1713593032
transform 1 0 1380 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1713593032
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _114_
timestamp 1713593032
transform -1 0 6256 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _115_
timestamp 1713593032
transform 1 0 1564 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _116_
timestamp 1713593032
transform -1 0 2760 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1713593032
transform 1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _118_
timestamp 1713593032
transform 1 0 5888 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _119_
timestamp 1713593032
transform -1 0 4692 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _120_
timestamp 1713593032
transform -1 0 5980 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1713593032
transform -1 0 6624 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _122_
timestamp 1713593032
transform 1 0 9476 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _123_
timestamp 1713593032
transform 1 0 9476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _124_
timestamp 1713593032
transform 1 0 4876 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1713593032
transform 1 0 5520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _126_
timestamp 1713593032
transform -1 0 3680 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _127_
timestamp 1713593032
transform -1 0 6532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _128_
timestamp 1713593032
transform -1 0 10396 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1713593032
transform 1 0 1472 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _130_
timestamp 1713593032
transform -1 0 2024 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _131_
timestamp 1713593032
transform 1 0 2852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _132_
timestamp 1713593032
transform 1 0 6808 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1713593032
transform 1 0 7820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _134_
timestamp 1713593032
transform -1 0 7912 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _135_
timestamp 1713593032
transform -1 0 5980 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _136_
timestamp 1713593032
transform -1 0 3312 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _137_
timestamp 1713593032
transform 1 0 4968 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1713593032
transform 1 0 7544 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _139_
timestamp 1713593032
transform -1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _140_
timestamp 1713593032
transform 1 0 3128 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2$2  _141_
timestamp 1713593032
transform -1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _142_
timestamp 1713593032
transform -1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _143_
timestamp 1713593032
transform -1 0 2484 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _144_
timestamp 1713593032
transform -1 0 5060 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _145_
timestamp 1713593032
transform 1 0 3864 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _146_
timestamp 1713593032
transform -1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _147_
timestamp 1713593032
transform 1 0 9660 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_2  _148_
timestamp 1713593032
transform -1 0 10488 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_2  _149_
timestamp 1713593032
transform -1 0 10304 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _150_
timestamp 1713593032
transform 1 0 4784 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _151_
timestamp 1713593032
transform -1 0 9844 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _152_
timestamp 1713593032
transform 1 0 2852 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1713593032
transform 1 0 4692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _154_
timestamp 1713593032
transform 1 0 2668 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _155_
timestamp 1713593032
transform -1 0 7176 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _156_
timestamp 1713593032
transform -1 0 10396 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1713593032
transform -1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _158_
timestamp 1713593032
transform -1 0 9660 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _159_
timestamp 1713593032
transform 1 0 2576 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _160_
timestamp 1713593032
transform -1 0 6900 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _161_
timestamp 1713593032
transform -1 0 8648 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1713593032
transform -1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _163_
timestamp 1713593032
transform -1 0 3588 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _164_
timestamp 1713593032
transform 1 0 2576 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _165_
timestamp 1713593032
transform -1 0 5796 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _166_
timestamp 1713593032
transform 1 0 2392 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _167_
timestamp 1713593032
transform -1 0 6164 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _168_
timestamp 1713593032
transform 1 0 2024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _169_
timestamp 1713593032
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _170_
timestamp 1713593032
transform -1 0 6900 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _171_
timestamp 1713593032
transform -1 0 9844 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _172_
timestamp 1713593032
transform 1 0 2668 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _173_
timestamp 1713593032
transform -1 0 9384 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _174_
timestamp 1713593032
transform -1 0 2576 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _175_
timestamp 1713593032
transform -1 0 5704 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _176_
timestamp 1713593032
transform -1 0 4324 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _177_
timestamp 1713593032
transform 1 0 4600 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1713593032
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _179_
timestamp 1713593032
transform 1 0 2392 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_2  _180_
timestamp 1713593032
transform 1 0 4692 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _181_
timestamp 1713593032
transform 1 0 4324 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1713593032
transform -1 0 8096 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2$2  _183_
timestamp 1713593032
transform -1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _184_
timestamp 1713593032
transform -1 0 7820 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _185_
timestamp 1713593032
transform -1 0 9476 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _186_
timestamp 1713593032
transform -1 0 7728 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1713593032
transform -1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _188_
timestamp 1713593032
transform -1 0 8832 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _189_
timestamp 1713593032
transform -1 0 2944 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _190_
timestamp 1713593032
transform 1 0 7084 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _191_
timestamp 1713593032
transform -1 0 5244 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _192_
timestamp 1713593032
transform -1 0 5336 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _193_
timestamp 1713593032
transform -1 0 9844 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _194_
timestamp 1713593032
transform 1 0 4692 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _195_
timestamp 1713593032
transform 1 0 1380 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _196_
timestamp 1713593032
transform -1 0 7820 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _197_
timestamp 1713593032
transform -1 0 5244 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _198_
timestamp 1713593032
transform -1 0 8004 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _199_
timestamp 1713593032
transform -1 0 5244 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _200_
timestamp 1713593032
transform 1 0 1380 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _201_
timestamp 1713593032
transform -1 0 4140 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _202_
timestamp 1713593032
transform 1 0 5980 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _203_
timestamp 1713593032
transform 1 0 6992 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _204_
timestamp 1713593032
transform 1 0 5612 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _205_
timestamp 1713593032
transform 1 0 6624 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _206_
timestamp 1713593032
transform 1 0 6532 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _207_
timestamp 1713593032
transform 1 0 8924 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _208_
timestamp 1713593032
transform 1 0 9016 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _209_
timestamp 1713593032
transform -1 0 9752 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _210_
timestamp 1713593032
transform 1 0 4324 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1713593032
transform -1 0 5336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1713593032
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1713593032
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1713593032
transform 1 0 5612 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1713593032
transform -1 0 5796 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1713593032
transform 1 0 7912 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_3
timestamp 1713593032
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_7
timestamp 1713593032
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18
timestamp 1713593032
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26
timestamp 1713593032
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1713593032
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_41
timestamp 1713593032
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_49
timestamp 1713593032
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1713593032
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1713593032
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1713593032
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1713593032
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1713593032
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_93
timestamp 1713593032
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_24
timestamp 1713593032
transform 1 0 3312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_52
timestamp 1713593032
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_61
timestamp 1713593032
transform 1 0 6716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_80
timestamp 1713593032
transform 1 0 8464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_88
timestamp 1713593032
transform 1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_3
timestamp 1713593032
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_12
timestamp 1713593032
transform 1 0 2208 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_23
timestamp 1713593032
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1713593032
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1713593032
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_37
timestamp 1713593032
transform 1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_65
timestamp 1713593032
transform 1 0 7084 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_72
timestamp 1713593032
transform 1 0 7728 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1713593032
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_90
timestamp 1713593032
transform 1 0 9384 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_96
timestamp 1713593032
transform 1 0 9936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_3
timestamp 1713593032
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_21
timestamp 1713593032
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_33
timestamp 1713593032
transform 1 0 4140 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_39
timestamp 1713593032
transform 1 0 4692 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_47
timestamp 1713593032
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1713593032
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_57
timestamp 1713593032
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_61
timestamp 1713593032
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_67
timestamp 1713593032
transform 1 0 7268 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_74
timestamp 1713593032
transform 1 0 7912 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_86
timestamp 1713593032
transform 1 0 9016 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_98
timestamp 1713593032
transform 1 0 10120 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1713593032
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_15
timestamp 1713593032
transform 1 0 2484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1713593032
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 1713593032
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_33
timestamp 1713593032
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_37
timestamp 1713593032
transform 1 0 4508 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_46
timestamp 1713593032
transform 1 0 5336 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_76
timestamp 1713593032
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1713593032
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_97
timestamp 1713593032
transform 1 0 10028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_10
timestamp 1713593032
transform 1 0 2024 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_16
timestamp 1713593032
transform 1 0 2576 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_22
timestamp 1713593032
transform 1 0 3128 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_28
timestamp 1713593032
transform 1 0 3680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_45
timestamp 1713593032
transform 1 0 5244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1713593032
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_57
timestamp 1713593032
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_94
timestamp 1713593032
transform 1 0 9752 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_101
timestamp 1713593032
transform 1 0 10396 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_20
timestamp 1713593032
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1713593032
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_37
timestamp 1713593032
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_42
timestamp 1713593032
transform 1 0 4968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_51
timestamp 1713593032
transform 1 0 5796 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_66
timestamp 1713593032
transform 1 0 7176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1713593032
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_94
timestamp 1713593032
transform 1 0 9752 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_98
timestamp 1713593032
transform 1 0 10120 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 1713593032
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_10
timestamp 1713593032
transform 1 0 2024 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_16
timestamp 1713593032
transform 1 0 2576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_51
timestamp 1713593032
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 1713593032
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_63
timestamp 1713593032
transform 1 0 6900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_98
timestamp 1713593032
transform 1 0 10120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 1713593032
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_20
timestamp 1713593032
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_45
timestamp 1713593032
transform 1 0 5244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_69
timestamp 1713593032
transform 1 0 7452 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_80
timestamp 1713593032
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_85
timestamp 1713593032
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_94
timestamp 1713593032
transform 1 0 9752 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_98
timestamp 1713593032
transform 1 0 10120 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_7
timestamp 1713593032
transform 1 0 1748 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_15
timestamp 1713593032
transform 1 0 2484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_33
timestamp 1713593032
transform 1 0 4140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1713593032
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_60
timestamp 1713593032
transform 1 0 6624 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_72
timestamp 1713593032
transform 1 0 7728 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_101
timestamp 1713593032
transform 1 0 10396 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1713593032
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1713593032
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1713593032
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 1713593032
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1713593032
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1713593032
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1713593032
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1713593032
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_85
timestamp 1713593032
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_93
timestamp 1713593032
transform 1 0 9660 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_20
timestamp 1713593032
transform 1 0 2944 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_32
timestamp 1713593032
transform 1 0 4048 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_43
timestamp 1713593032
transform 1 0 5060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_47
timestamp 1713593032
transform 1 0 5428 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1713593032
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1713593032
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1713593032
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_69
timestamp 1713593032
transform 1 0 7452 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_77
timestamp 1713593032
transform 1 0 8188 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_100
timestamp 1713593032
transform 1 0 10304 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1713593032
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_15
timestamp 1713593032
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_22
timestamp 1713593032
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 1713593032
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_39
timestamp 1713593032
transform 1 0 4692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_51
timestamp 1713593032
transform 1 0 5796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_76
timestamp 1713593032
transform 1 0 8096 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 1713593032
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_85
timestamp 1713593032
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_100
timestamp 1713593032
transform 1 0 10304 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_3
timestamp 1713593032
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_7
timestamp 1713593032
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_11
timestamp 1713593032
transform 1 0 2116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_16
timestamp 1713593032
transform 1 0 2576 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_26
timestamp 1713593032
transform 1 0 3496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_45
timestamp 1713593032
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_73
timestamp 1713593032
transform 1 0 7820 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_82
timestamp 1713593032
transform 1 0 8648 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_95
timestamp 1713593032
transform 1 0 9844 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1713593032
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_7
timestamp 1713593032
transform 1 0 1748 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_15
timestamp 1713593032
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_43
timestamp 1713593032
transform 1 0 5060 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_51
timestamp 1713593032
transform 1 0 5796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_75
timestamp 1713593032
transform 1 0 8004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_79
timestamp 1713593032
transform 1 0 8372 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1713593032
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_85
timestamp 1713593032
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_90
timestamp 1713593032
transform 1 0 9384 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_100
timestamp 1713593032
transform 1 0 10304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_3
timestamp 1713593032
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_12
timestamp 1713593032
transform 1 0 2208 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_18
timestamp 1713593032
transform 1 0 2760 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_22
timestamp 1713593032
transform 1 0 3128 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_34
timestamp 1713593032
transform 1 0 4232 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_46
timestamp 1713593032
transform 1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1713593032
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1713593032
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_76
timestamp 1713593032
transform 1 0 8096 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_7
timestamp 1713593032
transform 1 0 1748 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_13
timestamp 1713593032
transform 1 0 2300 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1713593032
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_29
timestamp 1713593032
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_39
timestamp 1713593032
transform 1 0 4692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_43
timestamp 1713593032
transform 1 0 5060 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_46
timestamp 1713593032
transform 1 0 5336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_53
timestamp 1713593032
transform 1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_57
timestamp 1713593032
transform 1 0 6348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_69
timestamp 1713593032
transform 1 0 7452 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_77
timestamp 1713593032
transform 1 0 8188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1713593032
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1713593032
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output3
timestamp 1713593032
transform 1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output4
timestamp 1713593032
transform -1 0 8556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 1713593032
transform 1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output6
timestamp 1713593032
transform 1 0 10212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output7
timestamp 1713593032
transform 1 0 10212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output8
timestamp 1713593032
transform 1 0 10212 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output9
timestamp 1713593032
transform 1 0 10212 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output10
timestamp 1713593032
transform 1 0 10212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output11
timestamp 1713593032
transform 1 0 10212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output12
timestamp 1713593032
transform 1 0 9936 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output13
timestamp 1713593032
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output14
timestamp 1713593032
transform 1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_17
timestamp 1713593032
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1713593032
transform -1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_18
timestamp 1713593032
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1713593032
transform -1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_19
timestamp 1713593032
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1713593032
transform -1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_20
timestamp 1713593032
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1713593032
transform -1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_21
timestamp 1713593032
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1713593032
transform -1 0 10764 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_22
timestamp 1713593032
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1713593032
transform -1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_23
timestamp 1713593032
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1713593032
transform -1 0 10764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_24
timestamp 1713593032
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1713593032
transform -1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_25
timestamp 1713593032
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1713593032
transform -1 0 10764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_26
timestamp 1713593032
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1713593032
transform -1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_27
timestamp 1713593032
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1713593032
transform -1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_28
timestamp 1713593032
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1713593032
transform -1 0 10764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_29
timestamp 1713593032
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1713593032
transform -1 0 10764 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_30
timestamp 1713593032
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1713593032
transform -1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_31
timestamp 1713593032
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1713593032
transform -1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_32
timestamp 1713593032
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1713593032
transform -1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_33
timestamp 1713593032
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1713593032
transform -1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_0_34
timestamp 1713593032
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_0_35
timestamp 1713593032
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_0_36
timestamp 1713593032
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_1_37
timestamp 1713593032
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_2_38
timestamp 1713593032
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_2_39
timestamp 1713593032
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_3_40
timestamp 1713593032
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_4_41
timestamp 1713593032
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_4_42
timestamp 1713593032
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_5_43
timestamp 1713593032
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_6_44
timestamp 1713593032
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_6_45
timestamp 1713593032
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_7_46
timestamp 1713593032
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_8_47
timestamp 1713593032
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_8_48
timestamp 1713593032
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_9_49
timestamp 1713593032
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_10_50
timestamp 1713593032
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_10_51
timestamp 1713593032
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_11_52
timestamp 1713593032
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_12_53
timestamp 1713593032
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_12_54
timestamp 1713593032
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_13_55
timestamp 1713593032
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_14_56
timestamp 1713593032
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_14_57
timestamp 1713593032
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_15_58
timestamp 1713593032
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_16_59
timestamp 1713593032
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_16_60
timestamp 1713593032
transform 1 0 6256 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1$3  TAP_TAPCELL_ROW_16_61
timestamp 1713593032
transform 1 0 8832 0 1 10880
box -38 -48 130 592
<< labels >>
rlabel metal1 s 5934 10880 5934 10880 4 VGND
rlabel metal1 s 5934 11424 5934 11424 4 VPWR
rlabel metal1 s 8468 5610 8468 5610 4 _000_
rlabel metal1 s 6854 4794 6854 4794 4 _002_
rlabel metal1 s 5167 6698 5167 6698 4 _003_
rlabel metal1 s 8050 5168 8050 5168 4 _004_
rlabel metal1 s 5285 7446 5285 7446 4 _006_
rlabel metal1 s 7774 9146 7774 9146 4 _008_
rlabel metal1 s 7134 5202 7134 5202 4 _010_
rlabel metal1 s 4462 5882 4462 5882 4 _013_
rlabel metal1 s 1794 6426 1794 6426 4 _014_
rlabel metal1 s 7212 3026 7212 3026 4 _015_
rlabel metal1 s 5832 3502 5832 3502 4 _016_
rlabel metal1 s 2530 2584 2530 2584 4 _017_
rlabel metal1 s 7038 7514 7038 7514 4 _019_
rlabel metal1 s 8678 10710 8678 10710 4 _020_
rlabel metal1 s 4687 3094 4687 3094 4 _022_
rlabel metal1 s 9568 3638 9568 3638 4 _024_
rlabel metal1 s 8556 10030 8556 10030 4 _025_
rlabel metal1 s 9660 9894 9660 9894 4 _026_
rlabel metal1 s 4692 4046 4692 4046 4 _027_
rlabel metal1 s 4692 5678 4692 5678 4 _029_
rlabel metal1 s 10166 5032 10166 5032 4 _030_
rlabel metal1 s 9246 6120 9246 6120 4 _033_
rlabel metal1 s 4738 10166 4738 10166 4 _034_
rlabel metal1 s 6854 5576 6854 5576 4 _035_
rlabel metal1 s 3312 3502 3312 3502 4 _036_
rlabel metal1 s 5972 5338 5972 5338 4 _037_
rlabel metal1 s 3634 4794 3634 4794 4 _038_
rlabel metal1 s 2714 2380 2714 2380 4 _039_
rlabel metal1 s 3634 9894 3634 9894 4 _040_
rlabel metal1 s 2438 2414 2438 2414 4 _041_
rlabel metal1 s 5658 5168 5658 5168 4 _043_
rlabel metal1 s 5014 9146 5014 9146 4 _044_
rlabel metal1 s 4562 8602 4562 8602 4 _047_
rlabel metal1 s 6394 7446 6394 7446 4 _048_
rlabel metal1 s 2530 6630 2530 6630 4 _049_
rlabel metal1 s 6302 10234 6302 10234 4 _051_
rlabel metal1 s 9154 5610 9154 5610 4 _053_
rlabel metal1 s 10258 8908 10258 8908 4 _055_
rlabel metal1 s 3680 6630 3680 6630 4 _057_
rlabel metal1 s 5888 2550 5888 2550 4 _059_
rlabel metal1 s 2714 10744 2714 10744 4 _060_
rlabel metal1 s 8234 8976 8234 8976 4 _061_
rlabel metal1 s 2116 6426 2116 6426 4 _062_
rlabel metal1 s 9509 8602 9509 8602 4 _063_
rlabel metal1 s 9798 5678 9798 5678 4 _064_
rlabel metal1 s 2898 6120 2898 6120 4 _065_
rlabel metal1 s 6118 4624 6118 4624 4 _067_
rlabel metal1 s 1840 5202 1840 5202 4 _068_
rlabel metal1 s 1702 4998 1702 4998 4 _069_
rlabel metal1 s 2645 10438 2645 10438 4 _071_
rlabel metal1 s 1886 3978 1886 3978 4 _072_
rlabel metal1 s 6118 10030 6118 10030 4 _074_
rlabel metal1 s 5474 7786 5474 7786 4 _075_
rlabel metal1 s 6394 4556 6394 4556 4 _076_
rlabel metal1 s 5244 4794 5244 4794 4 _079_
rlabel metal1 s 8694 7446 8694 7446 4 _081_
rlabel metal1 s 7222 4046 7222 4046 4 _085_
rlabel metal1 s 7314 3910 7314 3910 4 _086_
rlabel metal1 s 4784 2346 4784 2346 4 _088_
rlabel metal1 s 6900 2278 6900 2278 4 _089_
rlabel metal1 s 4324 4794 4324 4794 4 _090_
rlabel metal1 s 2024 2482 2024 2482 4 _091_
rlabel metal1 s 1702 2618 1702 2618 4 _093_
rlabel metal1 s 6900 6970 6900 6970 4 clknet_0_clk
rlabel metal1 s 1426 8500 1426 8500 4 clknet_1_0__leaf_clk
rlabel metal1 s 9706 5236 9706 5236 4 clknet_1_1__leaf_clk
rlabel metal1 s 8648 10642 8648 10642 4 counter\[0\]
rlabel metal1 s 4876 4590 4876 4590 4 counter\[10\]
rlabel metal1 s 6164 6358 6164 6358 4 counter\[2\]
rlabel metal1 s 3358 11118 3358 11118 4 counter\[3\]
rlabel metal1 s 2622 7990 2622 7990 4 counter\[4\]
rlabel metal1 s 7176 8602 7176 8602 4 counter\[5\]
rlabel metal1 s 6394 7242 6394 7242 4 counter\[6\]
rlabel metal1 s 6302 10064 6302 10064 4 counter\[7\]
rlabel metal1 s 1794 6868 1794 6868 4 counter\[8\]
rlabel metal1 s 2438 2482 2438 2482 4 net1
rlabel metal1 s 6670 6324 6670 6324 4 net10
rlabel metal1 s 7958 9928 7958 9928 4 net11
rlabel metal1 s 10028 9554 10028 9554 4 net12
rlabel metal1 s 7682 10778 7682 10778 4 net13
rlabel metal1 s 8326 11152 8326 11152 4 net14
rlabel metal1 s 1380 2414 1380 2414 4 net2
rlabel metal1 s 1932 2346 1932 2346 4 net3
rlabel metal1 s 5336 4046 5336 4046 4 net6
rlabel metal1 s 2898 5236 2898 5236 4 net7
rlabel metal1 s 10258 5712 10258 5712 4 net8
rlabel metal1 s 10258 6256 10258 6256 4 net9
rlabel metal1 s 10672 2278 10672 2278 4 ones[0]
rlabel metal1 s 9062 10778 9062 10778 4 ones[10]
flabel metal4 s 7604 2128 7924 11472 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2604 2128 2924 11472 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 6944 2128 7264 11472 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1944 2128 2264 11472 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
rlabel metal2 s 2622 5729 2622 5729 4 _001_
rlabel metal2 s 6578 4352 6578 4352 4 _005_
rlabel metal2 s 1697 3026 1697 3026 4 _007_
rlabel metal2 s 4926 5202 4926 5202 4 _009_
rlabel metal2 s 4926 9622 4926 9622 4 _011_
rlabel metal2 s 1150 6205 1150 6205 4 _012_
rlabel metal2 s 4738 9826 4738 9826 4 _018_
rlabel metal2 s 9434 5202 9434 5202 4 _021_
rlabel metal2 s 5014 3638 5014 3638 4 _023_
rlabel metal2 s 2530 6987 2530 6987 4 _028_
rlabel metal2 s 6946 5304 6946 5304 4 _031_
rlabel metal2 s 1334 5491 1334 5491 4 _032_
rlabel metal2 s 6486 8432 6486 8432 4 _042_
rlabel metal2 s 2346 9503 2346 9503 4 _045_
rlabel metal2 s 5566 5610 5566 5610 4 _046_
rlabel metal2 s 4830 4743 4830 4743 4 _050_
rlabel metal2 s 736 2074 736 2074 4 _054_
rlabel metal2 s 1886 10013 1886 10013 4 _056_
rlabel metal2 s 10074 4505 10074 4505 4 _058_
rlabel metal2 s 6946 7531 6946 7531 4 _066_
rlabel metal2 s 1978 5287 1978 5287 4 _070_
rlabel metal2 s 2346 10217 2346 10217 4 _073_
rlabel metal2 s 9890 4114 9890 4114 4 _077_
rlabel metal2 s 5114 4522 5114 4522 4 _078_
rlabel metal2 s 1978 6817 1978 6817 4 _080_
rlabel metal2 s 1702 10285 1702 10285 4 _082_
rlabel metal2 s 1886 5168 1886 5168 4 _083_
rlabel metal2 s 3542 8364 3542 8364 4 _084_
rlabel metal2 s 1242 6596 1242 6596 4 _092_
rlabel metal2 s 4646 10880 4646 10880 4 counter\[1\]
rlabel metal2 s 3266 6766 3266 6766 4 counter\[9\]
rlabel metal2 s 8326 10268 8326 10268 4 net4
rlabel metal2 s 9982 2587 9982 2587 4 net5
rlabel metal2 s 10166 2125 10166 2125 4 ones[1]
rlabel metal2 s 10442 3213 10442 3213 4 ones[2]
rlabel metal2 s 10442 4301 10442 4301 4 ones[3]
rlabel metal2 s 10442 5389 10442 5389 4 ones[4]
rlabel metal2 s 10442 6477 10442 6477 4 ones[5]
rlabel metal2 s 10442 7565 10442 7565 4 ones[6]
rlabel metal2 s 10442 8925 10442 8925 4 ones[7]
rlabel metal2 s 10166 9469 10166 9469 4 ones[8]
rlabel metal2 s 8786 10965 8786 10965 4 ones[9]
rlabel metal3 s 2070 3587 2070 3587 4 _052_
rlabel metal3 s 5037 9724 5037 9724 4 _087_
rlabel metal3 s 866 2244 866 2244 4 clk
rlabel metal3 s 0 11432 800 11552 4 pulse
port 15 nsew
rlabel metal3 s 9898 12852 9898 12852 4 ready
rlabel metal3 s 1096 6868 1096 6868 4 rst
flabel metal3 s 0 2184 800 2304 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 11108 824 11908 944 0 FreeSans 600 0 0 0 ones[0]
port 4 nsew
flabel metal3 s 11108 11704 11908 11824 0 FreeSans 600 0 0 0 ones[10]
port 5 nsew
flabel metal3 s 11108 1912 11908 2032 0 FreeSans 600 0 0 0 ones[1]
port 6 nsew
flabel metal3 s 11108 3000 11908 3120 0 FreeSans 600 0 0 0 ones[2]
port 7 nsew
flabel metal3 s 11108 4088 11908 4208 0 FreeSans 600 0 0 0 ones[3]
port 8 nsew
flabel metal3 s 11108 5176 11908 5296 0 FreeSans 600 0 0 0 ones[4]
port 9 nsew
flabel metal3 s 11108 6264 11908 6384 0 FreeSans 600 0 0 0 ones[5]
port 10 nsew
flabel metal3 s 11108 7352 11908 7472 0 FreeSans 600 0 0 0 ones[6]
port 11 nsew
flabel metal3 s 11108 8440 11908 8560 0 FreeSans 600 0 0 0 ones[7]
port 12 nsew
flabel metal3 s 11108 9528 11908 9648 0 FreeSans 600 0 0 0 ones[8]
port 13 nsew
flabel metal3 s 11108 10616 11908 10736 0 FreeSans 600 0 0 0 ones[9]
port 14 nsew
flabel metal3 s 400 11492 400 11492 0 FreeSans 600 0 0 0 pulse
flabel metal3 s 11108 12792 11908 12912 0 FreeSans 600 0 0 0 ready
port 16 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 rst
port 17 nsew
flabel metal5 s 1056 8676 10812 8996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3676 10812 3996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 8016 10812 8336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3016 10812 3336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 11908 14052
<< end >>
